* File: rcx_out.net
* Created: Tue Mar 26 09:42:55 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:42:55 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt NOR2X2  A B VDD VSS Y
* 
XM2/X1 Y B net010 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=2
XM1/X1 net010 A VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=2
XM3/X1 Y B VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM0/X1 Y A VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
*
* 
* .include "rcx_out.net.NOR2X2.pxi"
* BEGIN of "./rcx_out.net.NOR2X2.pxi"
* File: rcx_out.net.NOR2X2.pxi
* Created: Tue Mar 26 09:42:55 2019
* 

* END of "./rcx_out.net.NOR2X2.pxi"
* 
*
.ends
*
*

