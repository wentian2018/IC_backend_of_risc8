
module PCI_FIFO_1_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   g_array_0__4_, g_array_0__2_, g_array_1__5_, g_array_1__4_,
         g_array_1__2_, g_array_1__0_, g_array_2__5_, g_array_2__4_,
         g_array_2__3_, g_array_2__2_, g_array_2__1_, g_array_2__0_,
         g_array_3__5_, g_array_3__4_, g_array_3__3_, g_array_3__1_,
         pog_array_0__4_, pog_array_0__2_, pog_array_1__5_, pog_array_1__2_,
         pog_array_2__5_, pog_array_2__4_, pog_array_2__3_, pog_array_2__1_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  oai21d1 U1_4_2_5 ( .B1(pog_array_2__5_), .B2(g_array_2__2_), .A(
        g_array_2__5_), .ZN(g_array_3__5_) );
  oai21d1 U1_4_2_4 ( .B1(pog_array_2__4_), .B2(g_array_2__2_), .A(
        g_array_2__4_), .ZN(g_array_3__4_) );
  oai21d1 U1_4_2_3 ( .B1(pog_array_2__3_), .B2(g_array_2__2_), .A(
        g_array_2__3_), .ZN(g_array_3__3_) );
  oai21d1 U1_4_2_1 ( .B1(pog_array_2__1_), .B2(g_array_2__0_), .A(
        g_array_2__1_), .ZN(g_array_3__1_) );
  aoi21d1 U1_4_1_5 ( .B1(pog_array_1__5_), .B2(g_array_1__4_), .A(
        g_array_1__5_), .ZN(g_array_2__5_) );
  aoi21d1 U1_4_1_2 ( .B1(pog_array_1__2_), .B2(g_array_1__0_), .A(
        g_array_1__2_), .ZN(g_array_2__2_) );
  oai21d1 U1_4_0_4 ( .B1(pog_array_0__4_), .B2(g_array_2__3_), .A(
        g_array_0__4_), .ZN(g_array_1__4_) );
  oai21d1 U1_4_0_2 ( .B1(pog_array_0__2_), .B2(g_array_2__1_), .A(
        g_array_0__2_), .ZN(g_array_1__2_) );
  nd12d0 U1 ( .A1(pog_array_2__4_), .A2(pog_array_1__5_), .ZN(pog_array_2__5_)
         );
  nd02d0 U2 ( .A1(n1), .A2(n2), .ZN(pog_array_2__4_) );
  nr02d0 U3 ( .A1(pog_array_2__1_), .A2(pog_array_0__2_), .ZN(pog_array_1__2_)
         );
  inv0d0 U4 ( .I(n3), .ZN(pog_array_0__2_) );
  inv0d0 U5 ( .I(g_array_1__4_), .ZN(g_array_2__4_) );
  inv0d0 U6 ( .I(n4), .ZN(DIFF[6]) );
  xr03d1 U7 ( .A1(g_array_3__5_), .A2(B[6]), .A3(A[6]), .Z(n4) );
  mx02d0 U8 ( .I0(n5), .I1(n6), .S(g_array_3__4_), .Z(DIFF[5]) );
  nd12d0 U9 ( .A1(g_array_1__5_), .A2(pog_array_1__5_), .ZN(n6) );
  nd02d0 U10 ( .A1(B[5]), .A2(n7), .ZN(pog_array_1__5_) );
  nr02d0 U11 ( .A1(n7), .A2(B[5]), .ZN(g_array_1__5_) );
  inv0d0 U12 ( .I(A[5]), .ZN(n7) );
  xn02d1 U13 ( .A1(A[5]), .A2(B[5]), .ZN(n5) );
  mx02d0 U14 ( .I0(n8), .I1(n9), .S(g_array_3__3_), .Z(DIFF[4]) );
  nd02d0 U15 ( .A1(n1), .A2(g_array_0__4_), .ZN(n9) );
  nd02d0 U16 ( .A1(A[4]), .A2(n10), .ZN(g_array_0__4_) );
  inv0d0 U17 ( .I(pog_array_0__4_), .ZN(n1) );
  nr02d0 U18 ( .A1(n10), .A2(A[4]), .ZN(pog_array_0__4_) );
  inv0d0 U19 ( .I(B[4]), .ZN(n10) );
  xn02d1 U20 ( .A1(A[4]), .A2(B[4]), .ZN(n8) );
  xr02d1 U21 ( .A1(n11), .A2(g_array_2__2_), .Z(DIFF[3]) );
  nd02d0 U22 ( .A1(g_array_2__3_), .A2(n2), .ZN(n11) );
  inv0d0 U23 ( .I(pog_array_2__3_), .ZN(n2) );
  nr02d0 U24 ( .A1(n12), .A2(A[3]), .ZN(pog_array_2__3_) );
  nd02d0 U25 ( .A1(A[3]), .A2(n12), .ZN(g_array_2__3_) );
  inv0d0 U26 ( .I(B[3]), .ZN(n12) );
  mx02d0 U27 ( .I0(n13), .I1(n14), .S(g_array_3__1_), .Z(DIFF[2]) );
  nd02d0 U28 ( .A1(g_array_0__2_), .A2(n3), .ZN(n14) );
  nd02d0 U29 ( .A1(B[2]), .A2(n15), .ZN(n3) );
  nd12d0 U30 ( .A1(B[2]), .A2(A[2]), .ZN(g_array_0__2_) );
  xr02d1 U31 ( .A1(n15), .A2(B[2]), .Z(n13) );
  inv0d0 U32 ( .I(A[2]), .ZN(n15) );
  xr02d1 U33 ( .A1(g_array_1__0_), .A2(n16), .Z(DIFF[1]) );
  an12d1 U34 ( .A2(g_array_2__1_), .A1(pog_array_2__1_), .Z(n16) );
  nr02d0 U35 ( .A1(n17), .A2(A[1]), .ZN(pog_array_2__1_) );
  nd02d0 U36 ( .A1(A[1]), .A2(n17), .ZN(g_array_2__1_) );
  inv0d0 U37 ( .I(B[1]), .ZN(n17) );
  inv0d0 U38 ( .I(g_array_2__0_), .ZN(g_array_1__0_) );
  aor21d1 U39 ( .B1(A[0]), .B2(n18), .A(g_array_2__0_), .Z(DIFF[0]) );
  nr02d0 U40 ( .A1(n18), .A2(A[0]), .ZN(g_array_2__0_) );
  inv0d0 U41 ( .I(B[0]), .ZN(n18) );
endmodule


module PCI_FIFO_1_DW_inc_1 ( carry_in, a, carry_out, sum );
  input [6:0] a;
  output [6:0] sum;
  input carry_in;
  output carry_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  xr02d1 U2 ( .A1(a[6]), .A2(n1), .Z(sum[6]) );
  an12d1 U3 ( .A2(a[5]), .A1(n2), .Z(n1) );
  xn02d1 U4 ( .A1(a[5]), .A2(n2), .ZN(sum[5]) );
  nd02d0 U5 ( .A1(a[4]), .A2(n3), .ZN(n2) );
  xr02d1 U6 ( .A1(a[4]), .A2(n3), .Z(sum[4]) );
  nr03d0 U7 ( .A1(n4), .A2(n5), .A3(n6), .ZN(n3) );
  inv0d0 U8 ( .I(a[3]), .ZN(n6) );
  xr02d1 U9 ( .A1(a[3]), .A2(n7), .Z(sum[3]) );
  nr02d0 U10 ( .A1(n5), .A2(n4), .ZN(n7) );
  inv0d0 U11 ( .I(a[2]), .ZN(n4) );
  xn02d1 U12 ( .A1(a[2]), .A2(n5), .ZN(sum[2]) );
  nd03d0 U13 ( .A1(a[1]), .A2(a[0]), .A3(carry_in), .ZN(n5) );
  xn02d1 U14 ( .A1(a[1]), .A2(n8), .ZN(sum[1]) );
  nd02d0 U15 ( .A1(carry_in), .A2(a[0]), .ZN(n8) );
  xr02d1 U16 ( .A1(carry_in), .A2(a[0]), .Z(sum[0]) );
endmodule


module PCI_FIFO_1_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   g_array_0__4_, g_array_0__2_, g_array_1__5_, g_array_1__4_,
         g_array_1__2_, g_array_1__0_, g_array_2__5_, g_array_2__4_,
         g_array_2__3_, g_array_2__2_, g_array_2__1_, g_array_2__0_,
         g_array_3__5_, g_array_3__4_, g_array_3__3_, g_array_3__1_,
         pog_array_0__4_, pog_array_0__2_, pog_array_1__5_, pog_array_1__2_,
         pog_array_2__5_, pog_array_2__4_, pog_array_2__3_, pog_array_2__1_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  oai21d1 U1_4_2_5 ( .B1(pog_array_2__5_), .B2(g_array_2__2_), .A(
        g_array_2__5_), .ZN(g_array_3__5_) );
  oai21d1 U1_4_2_4 ( .B1(pog_array_2__4_), .B2(g_array_2__2_), .A(
        g_array_2__4_), .ZN(g_array_3__4_) );
  oai21d1 U1_4_2_3 ( .B1(pog_array_2__3_), .B2(g_array_2__2_), .A(
        g_array_2__3_), .ZN(g_array_3__3_) );
  oai21d1 U1_4_2_1 ( .B1(pog_array_2__1_), .B2(g_array_2__0_), .A(
        g_array_2__1_), .ZN(g_array_3__1_) );
  aoi21d1 U1_4_1_5 ( .B1(pog_array_1__5_), .B2(g_array_1__4_), .A(
        g_array_1__5_), .ZN(g_array_2__5_) );
  aoi21d1 U1_4_1_2 ( .B1(pog_array_1__2_), .B2(g_array_1__0_), .A(
        g_array_1__2_), .ZN(g_array_2__2_) );
  oai21d1 U1_4_0_4 ( .B1(pog_array_0__4_), .B2(g_array_2__3_), .A(
        g_array_0__4_), .ZN(g_array_1__4_) );
  oai21d1 U1_4_0_2 ( .B1(pog_array_0__2_), .B2(g_array_2__1_), .A(
        g_array_0__2_), .ZN(g_array_1__2_) );
  nd12d0 U1 ( .A1(pog_array_2__4_), .A2(pog_array_1__5_), .ZN(pog_array_2__5_)
         );
  nd02d0 U2 ( .A1(n1), .A2(n2), .ZN(pog_array_2__4_) );
  nr02d0 U3 ( .A1(pog_array_2__1_), .A2(pog_array_0__2_), .ZN(pog_array_1__2_)
         );
  inv0d0 U4 ( .I(n3), .ZN(pog_array_0__2_) );
  inv0d0 U5 ( .I(g_array_1__4_), .ZN(g_array_2__4_) );
  inv0d0 U6 ( .I(n4), .ZN(DIFF[6]) );
  xr03d1 U7 ( .A1(g_array_3__5_), .A2(B[6]), .A3(A[6]), .Z(n4) );
  mx02d0 U8 ( .I0(n5), .I1(n6), .S(g_array_3__4_), .Z(DIFF[5]) );
  nd12d0 U9 ( .A1(g_array_1__5_), .A2(pog_array_1__5_), .ZN(n6) );
  nd02d0 U10 ( .A1(B[5]), .A2(n7), .ZN(pog_array_1__5_) );
  nr02d0 U11 ( .A1(n7), .A2(B[5]), .ZN(g_array_1__5_) );
  inv0d0 U12 ( .I(A[5]), .ZN(n7) );
  xn02d1 U13 ( .A1(A[5]), .A2(B[5]), .ZN(n5) );
  mx02d0 U14 ( .I0(n8), .I1(n9), .S(g_array_3__3_), .Z(DIFF[4]) );
  nd02d0 U15 ( .A1(n1), .A2(g_array_0__4_), .ZN(n9) );
  nd02d0 U16 ( .A1(A[4]), .A2(n10), .ZN(g_array_0__4_) );
  inv0d0 U17 ( .I(pog_array_0__4_), .ZN(n1) );
  nr02d0 U18 ( .A1(n10), .A2(A[4]), .ZN(pog_array_0__4_) );
  inv0d0 U19 ( .I(B[4]), .ZN(n10) );
  xn02d1 U20 ( .A1(A[4]), .A2(B[4]), .ZN(n8) );
  xr02d1 U21 ( .A1(n11), .A2(g_array_2__2_), .Z(DIFF[3]) );
  nd02d0 U22 ( .A1(g_array_2__3_), .A2(n2), .ZN(n11) );
  inv0d0 U23 ( .I(pog_array_2__3_), .ZN(n2) );
  nr02d0 U24 ( .A1(n12), .A2(A[3]), .ZN(pog_array_2__3_) );
  nd02d0 U25 ( .A1(A[3]), .A2(n12), .ZN(g_array_2__3_) );
  inv0d0 U26 ( .I(B[3]), .ZN(n12) );
  mx02d0 U27 ( .I0(n13), .I1(n14), .S(g_array_3__1_), .Z(DIFF[2]) );
  nd02d0 U28 ( .A1(g_array_0__2_), .A2(n3), .ZN(n14) );
  nd02d0 U29 ( .A1(B[2]), .A2(n15), .ZN(n3) );
  nd12d0 U30 ( .A1(B[2]), .A2(A[2]), .ZN(g_array_0__2_) );
  xr02d1 U31 ( .A1(n15), .A2(B[2]), .Z(n13) );
  inv0d0 U32 ( .I(A[2]), .ZN(n15) );
  xr02d1 U33 ( .A1(g_array_1__0_), .A2(n16), .Z(DIFF[1]) );
  an12d1 U34 ( .A2(g_array_2__1_), .A1(pog_array_2__1_), .Z(n16) );
  nr02d0 U35 ( .A1(n17), .A2(A[1]), .ZN(pog_array_2__1_) );
  nd02d0 U36 ( .A1(A[1]), .A2(n17), .ZN(g_array_2__1_) );
  inv0d0 U37 ( .I(B[1]), .ZN(n17) );
  inv0d0 U38 ( .I(g_array_2__0_), .ZN(g_array_1__0_) );
  aor21d1 U39 ( .B1(A[0]), .B2(n18), .A(g_array_2__0_), .Z(DIFF[0]) );
  nr02d0 U40 ( .A1(n18), .A2(A[0]), .ZN(g_array_2__0_) );
  inv0d0 U41 ( .I(B[0]), .ZN(n18) );
endmodule


module PCI_FIFO_1_DW_inc_0 ( carry_in, a, carry_out, sum );
  input [6:0] a;
  output [6:0] sum;
  input carry_in;
  output carry_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  xr02d1 U2 ( .A1(a[6]), .A2(n1), .Z(sum[6]) );
  an12d1 U3 ( .A2(a[5]), .A1(n2), .Z(n1) );
  xn02d1 U4 ( .A1(a[5]), .A2(n2), .ZN(sum[5]) );
  nd02d0 U5 ( .A1(a[4]), .A2(n3), .ZN(n2) );
  xr02d1 U6 ( .A1(a[4]), .A2(n3), .Z(sum[4]) );
  nr03d0 U7 ( .A1(n4), .A2(n5), .A3(n6), .ZN(n3) );
  inv0d0 U8 ( .I(a[3]), .ZN(n6) );
  xr02d1 U9 ( .A1(a[3]), .A2(n7), .Z(sum[3]) );
  nr02d0 U10 ( .A1(n5), .A2(n4), .ZN(n7) );
  inv0d0 U11 ( .I(a[2]), .ZN(n4) );
  xn02d1 U12 ( .A1(a[2]), .A2(n5), .ZN(sum[2]) );
  nd03d0 U13 ( .A1(a[1]), .A2(a[0]), .A3(carry_in), .ZN(n5) );
  xn02d1 U14 ( .A1(a[1]), .A2(n8), .ZN(sum[1]) );
  nd02d0 U15 ( .A1(carry_in), .A2(a[0]), .ZN(n8) );
  xr02d1 U16 ( .A1(carry_in), .A2(a[0]), .Z(sum[0]) );
endmodule


module PCI_FIFO_0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   g_array_0__4_, g_array_0__2_, g_array_1__5_, g_array_1__4_,
         g_array_1__2_, g_array_1__0_, g_array_2__5_, g_array_2__4_,
         g_array_2__3_, g_array_2__2_, g_array_2__1_, g_array_2__0_,
         g_array_3__5_, g_array_3__4_, g_array_3__3_, g_array_3__1_,
         pog_array_0__4_, pog_array_0__2_, pog_array_1__5_, pog_array_1__2_,
         pog_array_2__5_, pog_array_2__4_, pog_array_2__3_, pog_array_2__1_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  oai21d1 U1_4_2_5 ( .B1(pog_array_2__5_), .B2(g_array_2__2_), .A(
        g_array_2__5_), .ZN(g_array_3__5_) );
  oai21d1 U1_4_2_4 ( .B1(pog_array_2__4_), .B2(g_array_2__2_), .A(
        g_array_2__4_), .ZN(g_array_3__4_) );
  oai21d1 U1_4_2_3 ( .B1(pog_array_2__3_), .B2(g_array_2__2_), .A(
        g_array_2__3_), .ZN(g_array_3__3_) );
  oai21d1 U1_4_2_1 ( .B1(pog_array_2__1_), .B2(g_array_2__0_), .A(
        g_array_2__1_), .ZN(g_array_3__1_) );
  aoi21d1 U1_4_1_5 ( .B1(pog_array_1__5_), .B2(g_array_1__4_), .A(
        g_array_1__5_), .ZN(g_array_2__5_) );
  aoi21d1 U1_4_1_2 ( .B1(pog_array_1__2_), .B2(g_array_1__0_), .A(
        g_array_1__2_), .ZN(g_array_2__2_) );
  oai21d1 U1_4_0_4 ( .B1(pog_array_0__4_), .B2(g_array_2__3_), .A(
        g_array_0__4_), .ZN(g_array_1__4_) );
  oai21d1 U1_4_0_2 ( .B1(pog_array_0__2_), .B2(g_array_2__1_), .A(
        g_array_0__2_), .ZN(g_array_1__2_) );
  nd12d0 U1 ( .A1(pog_array_2__4_), .A2(pog_array_1__5_), .ZN(pog_array_2__5_)
         );
  nd02d0 U2 ( .A1(n1), .A2(n2), .ZN(pog_array_2__4_) );
  nr02d0 U3 ( .A1(pog_array_2__1_), .A2(pog_array_0__2_), .ZN(pog_array_1__2_)
         );
  inv0d0 U4 ( .I(n3), .ZN(pog_array_0__2_) );
  inv0d0 U5 ( .I(g_array_1__4_), .ZN(g_array_2__4_) );
  inv0d0 U6 ( .I(n4), .ZN(DIFF[6]) );
  xr03d1 U7 ( .A1(g_array_3__5_), .A2(B[6]), .A3(A[6]), .Z(n4) );
  mx02d0 U8 ( .I0(n5), .I1(n6), .S(g_array_3__4_), .Z(DIFF[5]) );
  nd12d0 U9 ( .A1(g_array_1__5_), .A2(pog_array_1__5_), .ZN(n6) );
  nd02d0 U10 ( .A1(B[5]), .A2(n7), .ZN(pog_array_1__5_) );
  nr02d0 U11 ( .A1(n7), .A2(B[5]), .ZN(g_array_1__5_) );
  inv0d0 U12 ( .I(A[5]), .ZN(n7) );
  xn02d1 U13 ( .A1(A[5]), .A2(B[5]), .ZN(n5) );
  mx02d0 U14 ( .I0(n8), .I1(n9), .S(g_array_3__3_), .Z(DIFF[4]) );
  nd02d0 U15 ( .A1(n1), .A2(g_array_0__4_), .ZN(n9) );
  nd02d0 U16 ( .A1(A[4]), .A2(n10), .ZN(g_array_0__4_) );
  inv0d0 U17 ( .I(pog_array_0__4_), .ZN(n1) );
  nr02d0 U18 ( .A1(n10), .A2(A[4]), .ZN(pog_array_0__4_) );
  inv0d0 U19 ( .I(B[4]), .ZN(n10) );
  xn02d1 U20 ( .A1(A[4]), .A2(B[4]), .ZN(n8) );
  xr02d1 U21 ( .A1(n11), .A2(g_array_2__2_), .Z(DIFF[3]) );
  nd02d0 U22 ( .A1(g_array_2__3_), .A2(n2), .ZN(n11) );
  inv0d0 U23 ( .I(pog_array_2__3_), .ZN(n2) );
  nr02d0 U24 ( .A1(n12), .A2(A[3]), .ZN(pog_array_2__3_) );
  nd02d0 U25 ( .A1(A[3]), .A2(n12), .ZN(g_array_2__3_) );
  inv0d0 U26 ( .I(B[3]), .ZN(n12) );
  mx02d0 U27 ( .I0(n13), .I1(n14), .S(g_array_3__1_), .Z(DIFF[2]) );
  nd02d0 U28 ( .A1(g_array_0__2_), .A2(n3), .ZN(n14) );
  nd02d0 U29 ( .A1(B[2]), .A2(n15), .ZN(n3) );
  nd12d0 U30 ( .A1(B[2]), .A2(A[2]), .ZN(g_array_0__2_) );
  xr02d1 U31 ( .A1(n15), .A2(B[2]), .Z(n13) );
  inv0d0 U32 ( .I(A[2]), .ZN(n15) );
  xr02d1 U33 ( .A1(g_array_1__0_), .A2(n16), .Z(DIFF[1]) );
  an12d1 U34 ( .A2(g_array_2__1_), .A1(pog_array_2__1_), .Z(n16) );
  nr02d0 U35 ( .A1(n17), .A2(A[1]), .ZN(pog_array_2__1_) );
  nd02d0 U36 ( .A1(A[1]), .A2(n17), .ZN(g_array_2__1_) );
  inv0d0 U37 ( .I(B[1]), .ZN(n17) );
  inv0d0 U38 ( .I(g_array_2__0_), .ZN(g_array_1__0_) );
  aor21d1 U39 ( .B1(A[0]), .B2(n18), .A(g_array_2__0_), .Z(DIFF[0]) );
  nr02d0 U40 ( .A1(n18), .A2(A[0]), .ZN(g_array_2__0_) );
  inv0d0 U41 ( .I(B[0]), .ZN(n18) );
endmodule


module PCI_FIFO_0_DW_inc_1 ( carry_in, a, carry_out, sum );
  input [6:0] a;
  output [6:0] sum;
  input carry_in;
  output carry_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  xr02d1 U2 ( .A1(a[6]), .A2(n1), .Z(sum[6]) );
  an12d1 U3 ( .A2(a[5]), .A1(n2), .Z(n1) );
  xn02d1 U4 ( .A1(a[5]), .A2(n2), .ZN(sum[5]) );
  nd02d0 U5 ( .A1(a[4]), .A2(n3), .ZN(n2) );
  xr02d1 U6 ( .A1(a[4]), .A2(n3), .Z(sum[4]) );
  nr03d0 U7 ( .A1(n4), .A2(n5), .A3(n6), .ZN(n3) );
  inv0d0 U8 ( .I(a[3]), .ZN(n6) );
  xr02d1 U9 ( .A1(a[3]), .A2(n7), .Z(sum[3]) );
  nr02d0 U10 ( .A1(n5), .A2(n4), .ZN(n7) );
  inv0d0 U11 ( .I(a[2]), .ZN(n4) );
  xn02d1 U12 ( .A1(a[2]), .A2(n5), .ZN(sum[2]) );
  nd03d0 U13 ( .A1(a[1]), .A2(a[0]), .A3(carry_in), .ZN(n5) );
  xn02d1 U14 ( .A1(a[1]), .A2(n8), .ZN(sum[1]) );
  nd02d0 U15 ( .A1(carry_in), .A2(a[0]), .ZN(n8) );
  xr02d1 U16 ( .A1(carry_in), .A2(a[0]), .Z(sum[0]) );
endmodule


module PCI_FIFO_0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   g_array_0__4_, g_array_0__2_, g_array_1__5_, g_array_1__4_,
         g_array_1__2_, g_array_1__0_, g_array_2__5_, g_array_2__4_,
         g_array_2__3_, g_array_2__2_, g_array_2__1_, g_array_2__0_,
         g_array_3__5_, g_array_3__4_, g_array_3__3_, g_array_3__1_,
         pog_array_0__4_, pog_array_0__2_, pog_array_1__5_, pog_array_1__2_,
         pog_array_2__5_, pog_array_2__4_, pog_array_2__3_, pog_array_2__1_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  oai21d1 U1_4_2_5 ( .B1(pog_array_2__5_), .B2(g_array_2__2_), .A(
        g_array_2__5_), .ZN(g_array_3__5_) );
  oai21d1 U1_4_2_4 ( .B1(pog_array_2__4_), .B2(g_array_2__2_), .A(
        g_array_2__4_), .ZN(g_array_3__4_) );
  oai21d1 U1_4_2_3 ( .B1(pog_array_2__3_), .B2(g_array_2__2_), .A(
        g_array_2__3_), .ZN(g_array_3__3_) );
  oai21d1 U1_4_2_1 ( .B1(pog_array_2__1_), .B2(g_array_2__0_), .A(
        g_array_2__1_), .ZN(g_array_3__1_) );
  aoi21d1 U1_4_1_5 ( .B1(pog_array_1__5_), .B2(g_array_1__4_), .A(
        g_array_1__5_), .ZN(g_array_2__5_) );
  aoi21d1 U1_4_1_2 ( .B1(pog_array_1__2_), .B2(g_array_1__0_), .A(
        g_array_1__2_), .ZN(g_array_2__2_) );
  oai21d1 U1_4_0_4 ( .B1(pog_array_0__4_), .B2(g_array_2__3_), .A(
        g_array_0__4_), .ZN(g_array_1__4_) );
  oai21d1 U1_4_0_2 ( .B1(pog_array_0__2_), .B2(g_array_2__1_), .A(
        g_array_0__2_), .ZN(g_array_1__2_) );
  nd12d0 U1 ( .A1(pog_array_2__4_), .A2(pog_array_1__5_), .ZN(pog_array_2__5_)
         );
  nd02d0 U2 ( .A1(n1), .A2(n2), .ZN(pog_array_2__4_) );
  nr02d0 U3 ( .A1(pog_array_2__1_), .A2(pog_array_0__2_), .ZN(pog_array_1__2_)
         );
  inv0d0 U4 ( .I(n3), .ZN(pog_array_0__2_) );
  inv0d0 U5 ( .I(g_array_1__4_), .ZN(g_array_2__4_) );
  inv0d0 U6 ( .I(n4), .ZN(DIFF[6]) );
  xr03d1 U7 ( .A1(g_array_3__5_), .A2(B[6]), .A3(A[6]), .Z(n4) );
  mx02d0 U8 ( .I0(n5), .I1(n6), .S(g_array_3__4_), .Z(DIFF[5]) );
  nd12d0 U9 ( .A1(g_array_1__5_), .A2(pog_array_1__5_), .ZN(n6) );
  nd02d0 U10 ( .A1(B[5]), .A2(n7), .ZN(pog_array_1__5_) );
  nr02d0 U11 ( .A1(n7), .A2(B[5]), .ZN(g_array_1__5_) );
  inv0d0 U12 ( .I(A[5]), .ZN(n7) );
  xn02d1 U13 ( .A1(A[5]), .A2(B[5]), .ZN(n5) );
  mx02d0 U14 ( .I0(n8), .I1(n9), .S(g_array_3__3_), .Z(DIFF[4]) );
  nd02d0 U15 ( .A1(n1), .A2(g_array_0__4_), .ZN(n9) );
  nd02d0 U16 ( .A1(A[4]), .A2(n10), .ZN(g_array_0__4_) );
  inv0d0 U17 ( .I(pog_array_0__4_), .ZN(n1) );
  nr02d0 U18 ( .A1(n10), .A2(A[4]), .ZN(pog_array_0__4_) );
  inv0d0 U19 ( .I(B[4]), .ZN(n10) );
  xn02d1 U20 ( .A1(A[4]), .A2(B[4]), .ZN(n8) );
  xr02d1 U21 ( .A1(n11), .A2(g_array_2__2_), .Z(DIFF[3]) );
  nd02d0 U22 ( .A1(g_array_2__3_), .A2(n2), .ZN(n11) );
  inv0d0 U23 ( .I(pog_array_2__3_), .ZN(n2) );
  nr02d0 U24 ( .A1(n12), .A2(A[3]), .ZN(pog_array_2__3_) );
  nd02d0 U25 ( .A1(A[3]), .A2(n12), .ZN(g_array_2__3_) );
  inv0d0 U26 ( .I(B[3]), .ZN(n12) );
  mx02d0 U27 ( .I0(n13), .I1(n14), .S(g_array_3__1_), .Z(DIFF[2]) );
  nd02d0 U28 ( .A1(g_array_0__2_), .A2(n3), .ZN(n14) );
  nd02d0 U29 ( .A1(B[2]), .A2(n15), .ZN(n3) );
  nd12d0 U30 ( .A1(B[2]), .A2(A[2]), .ZN(g_array_0__2_) );
  xr02d1 U31 ( .A1(n15), .A2(B[2]), .Z(n13) );
  inv0d0 U32 ( .I(A[2]), .ZN(n15) );
  xr02d1 U33 ( .A1(g_array_1__0_), .A2(n16), .Z(DIFF[1]) );
  an12d1 U34 ( .A2(g_array_2__1_), .A1(pog_array_2__1_), .Z(n16) );
  nr02d0 U35 ( .A1(n17), .A2(A[1]), .ZN(pog_array_2__1_) );
  nd02d0 U36 ( .A1(A[1]), .A2(n17), .ZN(g_array_2__1_) );
  inv0d0 U37 ( .I(B[1]), .ZN(n17) );
  inv0d0 U38 ( .I(g_array_2__0_), .ZN(g_array_1__0_) );
  aor21d1 U39 ( .B1(A[0]), .B2(n18), .A(g_array_2__0_), .Z(DIFF[0]) );
  nr02d0 U40 ( .A1(n18), .A2(A[0]), .ZN(g_array_2__0_) );
  inv0d0 U41 ( .I(B[0]), .ZN(n18) );
endmodule


module PCI_FIFO_0_DW_inc_0 ( carry_in, a, carry_out, sum );
  input [6:0] a;
  output [6:0] sum;
  input carry_in;
  output carry_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  xr02d1 U2 ( .A1(a[6]), .A2(n1), .Z(sum[6]) );
  an12d1 U3 ( .A2(a[5]), .A1(n2), .Z(n1) );
  xn02d1 U4 ( .A1(a[5]), .A2(n2), .ZN(sum[5]) );
  nd02d0 U5 ( .A1(a[4]), .A2(n3), .ZN(n2) );
  xr02d1 U6 ( .A1(a[4]), .A2(n3), .Z(sum[4]) );
  nr03d0 U7 ( .A1(n4), .A2(n5), .A3(n6), .ZN(n3) );
  inv0d0 U8 ( .I(a[3]), .ZN(n6) );
  xr02d1 U9 ( .A1(a[3]), .A2(n7), .Z(sum[3]) );
  nr02d0 U10 ( .A1(n5), .A2(n4), .ZN(n7) );
  inv0d0 U11 ( .I(a[2]), .ZN(n4) );
  xn02d1 U12 ( .A1(a[2]), .A2(n5), .ZN(sum[2]) );
  nd03d0 U13 ( .A1(a[1]), .A2(a[0]), .A3(carry_in), .ZN(n5) );
  xn02d1 U14 ( .A1(a[1]), .A2(n8), .ZN(sum[1]) );
  nd02d0 U15 ( .A1(carry_in), .A2(a[0]), .ZN(n8) );
  xr02d1 U16 ( .A1(carry_in), .A2(a[0]), .Z(sum[0]) );
endmodule


module SDRAM_FIFO_1_DW_FIFOCTL_IF_1 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [3:0] other_addr_g;
  output [3:0] word_count;
  output [2:0] this_addr;
  output [3:0] this_addr_g;
  output [3:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_3_, sync_2_, sync_1_, sync_0_, count_int_3_, empty_int, N6, N7,
         N8, N9, N10, N11, N12, N18, N19, N20, N21, N22, N23, n15, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50;

  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrn1 empty_int_reg ( .D(N18), .SD(count_int_3_), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(n15) );
  sdcrq1 count_int_reg_0_ ( .D(N6), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 count_int_reg_1_ ( .D(N7), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_2_ ( .D(N8), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_3_ ( .D(N9), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_int_3_) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N12), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N9), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N11), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N10), .SD(sync_3_), .SC(test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrq1 error_int_reg ( .D(N23), .SD(n15), .SC(test_se), .CP(clk), .CDN(rst_n), .Q(error) );
  sdcrn1 almost_empty_int_reg ( .D(N19), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrq1 half_full_int_reg ( .D(N20), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(N21), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrq1 full_int_reg ( .D(N22), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  inv0d1 U20 ( .I(n15), .ZN(empty_int) );
  aor21d1 U25 ( .B1(empty), .B2(n20), .A(error), .Z(N23) );
  inv0d0 U26 ( .I(empty_int), .ZN(empty) );
  nr04d0 U27 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(N22) );
  aor21d1 U28 ( .B1(n21), .B2(n22), .A(n25), .Z(N21) );
  inv0d0 U29 ( .I(n26), .ZN(n22) );
  aor21d1 U30 ( .B1(n21), .B2(n24), .A(N20), .Z(N19) );
  or03d0 U31 ( .A1(n21), .A2(N20), .A3(n24), .Z(N18) );
  xn02d1 U32 ( .A1(n27), .A2(n28), .ZN(n24) );
  nd02d0 U33 ( .A1(n23), .A2(n26), .ZN(N20) );
  xn02d1 U34 ( .A1(n29), .A2(n30), .ZN(n26) );
  an02d0 U35 ( .A1(n31), .A2(n32), .Z(n30) );
  nd02d0 U36 ( .A1(n33), .A2(n34), .ZN(n29) );
  inv0d0 U37 ( .I(n25), .ZN(n23) );
  xr03d1 U38 ( .A1(sync_3_), .A2(n35), .A3(n36), .Z(n25) );
  oai221d1 U39 ( .B1(n37), .B2(n31), .C1(n37), .C2(n32), .A(n34), .ZN(n35) );
  nd02d0 U40 ( .A1(n38), .A2(n39), .ZN(n34) );
  nd02d0 U41 ( .A1(n40), .A2(n41), .ZN(n32) );
  inv0d0 U42 ( .I(n33), .ZN(n37) );
  nd02d0 U43 ( .A1(n42), .A2(N8), .ZN(n33) );
  xn02d1 U44 ( .A1(n43), .A2(n40), .ZN(n21) );
  or02d0 U45 ( .A1(n28), .A2(n27), .Z(n40) );
  xn02d1 U46 ( .A1(n44), .A2(sync_0_), .ZN(n28) );
  nd02d0 U47 ( .A1(n31), .A2(n41), .ZN(n43) );
  nd02d0 U48 ( .A1(n44), .A2(N7), .ZN(n41) );
  inv0d0 U49 ( .I(n45), .ZN(n44) );
  nd02d0 U50 ( .A1(n45), .A2(n46), .ZN(n31) );
  xn02d1 U51 ( .A1(n42), .A2(sync_1_), .ZN(n45) );
  inv0d0 U52 ( .I(n38), .ZN(n42) );
  xr02d1 U53 ( .A1(sync_3_), .A2(sync_2_), .Z(n38) );
  xr02d1 U54 ( .A1(n36), .A2(n39), .Z(N12) );
  inv0d0 U55 ( .I(N9), .ZN(n36) );
  xn02d1 U56 ( .A1(n47), .A2(count_int_3_), .ZN(N9) );
  nd02d0 U57 ( .A1(this_addr[2]), .A2(n48), .ZN(n47) );
  xr02d1 U58 ( .A1(N8), .A2(N7), .Z(N11) );
  inv0d0 U59 ( .I(n46), .ZN(N7) );
  inv0d0 U60 ( .I(n39), .ZN(N8) );
  xn02d1 U61 ( .A1(this_addr[2]), .A2(n48), .ZN(n39) );
  an12d1 U62 ( .A2(this_addr[1]), .A1(n49), .Z(n48) );
  xn02d1 U63 ( .A1(n46), .A2(N6), .ZN(N10) );
  inv0d0 U64 ( .I(n27), .ZN(N6) );
  xr02d1 U65 ( .A1(n50), .A2(this_addr[0]), .Z(n27) );
  nd02d0 U66 ( .A1(empty_int), .A2(n20), .ZN(n50) );
  xr02d1 U67 ( .A1(n49), .A2(this_addr[1]), .Z(n46) );
  nd03d0 U68 ( .A1(empty_int), .A2(n20), .A3(this_addr[0]), .ZN(n49) );
  inv0d0 U69 ( .I(inc_req_n), .ZN(n20) );
endmodule


module SDRAM_FIFO_1_DW_FIFOCTL_IF_0 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [3:0] other_addr_g;
  output [3:0] word_count;
  output [2:0] this_addr;
  output [3:0] this_addr_g;
  output [3:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_3_, sync_2_, sync_1_, sync_0_, count_int_3_, N6, N7, N8, N9, N10,
         N11, N12, N18, N19, N20, N21, N22, N23, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48;

  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrq1 full_int_reg ( .D(N22), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  sdcrq1 count_int_reg_0_ ( .D(N6), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 count_int_reg_1_ ( .D(N7), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_2_ ( .D(N8), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_3_ ( .D(N9), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_int_3_) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N9), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N12), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N11), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 half_full_int_reg ( .D(N20), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(N21), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrn1 almost_empty_int_reg ( .D(N19), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrn1 empty_int_reg ( .D(N18), .SD(count_int_3_), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(empty) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N10), .SD(sync_3_), .SC(test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrq1 error_int_reg ( .D(N23), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  aor21d1 U24 ( .B1(full), .B2(n19), .A(error), .Z(N23) );
  inv0d0 U25 ( .I(inc_req_n), .ZN(n19) );
  nr04d0 U26 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(N22) );
  aor21d1 U27 ( .B1(n20), .B2(n21), .A(n24), .Z(N21) );
  inv0d0 U28 ( .I(n25), .ZN(n21) );
  aor21d1 U29 ( .B1(n20), .B2(n23), .A(N20), .Z(N19) );
  or03d0 U30 ( .A1(n20), .A2(N20), .A3(n23), .Z(N18) );
  xn02d1 U31 ( .A1(n26), .A2(n27), .ZN(n23) );
  nd02d0 U32 ( .A1(n22), .A2(n25), .ZN(N20) );
  xn02d1 U33 ( .A1(n28), .A2(n29), .ZN(n25) );
  an12d1 U34 ( .A2(n30), .A1(n31), .Z(n29) );
  nd02d0 U35 ( .A1(n32), .A2(n33), .ZN(n28) );
  inv0d0 U36 ( .I(n24), .ZN(n22) );
  xr03d1 U37 ( .A1(sync_3_), .A2(n34), .A3(n35), .Z(n24) );
  oai221d1 U38 ( .B1(n31), .B2(n33), .C1(n31), .C2(n32), .A(n30), .ZN(n34) );
  nd02d0 U39 ( .A1(n36), .A2(N8), .ZN(n30) );
  nd02d0 U40 ( .A1(n37), .A2(n38), .ZN(n32) );
  nr02d0 U41 ( .A1(n36), .A2(N8), .ZN(n31) );
  inv0d0 U42 ( .I(n39), .ZN(N8) );
  xr02d1 U43 ( .A1(n37), .A2(n40), .Z(n20) );
  an02d0 U44 ( .A1(n38), .A2(n33), .Z(n40) );
  nd02d0 U45 ( .A1(n41), .A2(N7), .ZN(n33) );
  nd02d0 U46 ( .A1(n42), .A2(n43), .ZN(n38) );
  nd02d0 U47 ( .A1(n27), .A2(n26), .ZN(n37) );
  xn02d1 U48 ( .A1(n41), .A2(sync_0_), .ZN(n27) );
  inv0d0 U49 ( .I(n42), .ZN(n41) );
  xn02d1 U50 ( .A1(n36), .A2(sync_1_), .ZN(n42) );
  xn02d1 U51 ( .A1(sync_3_), .A2(sync_2_), .ZN(n36) );
  xr02d1 U52 ( .A1(n35), .A2(n39), .Z(N12) );
  inv0d0 U53 ( .I(N9), .ZN(n35) );
  xn02d1 U54 ( .A1(n44), .A2(count_int_3_), .ZN(N9) );
  nd02d0 U55 ( .A1(this_addr[2]), .A2(n45), .ZN(n44) );
  xn02d1 U56 ( .A1(n39), .A2(N7), .ZN(N11) );
  inv0d0 U57 ( .I(n43), .ZN(N7) );
  xn02d1 U58 ( .A1(this_addr[2]), .A2(n45), .ZN(n39) );
  an02d0 U59 ( .A1(this_addr[1]), .A2(n46), .Z(n45) );
  xr02d1 U60 ( .A1(n43), .A2(n26), .Z(N10) );
  inv0d0 U61 ( .I(N6), .ZN(n26) );
  xn02d1 U62 ( .A1(n47), .A2(n48), .ZN(N6) );
  nr02d0 U63 ( .A1(full), .A2(inc_req_n), .ZN(n48) );
  xn02d1 U64 ( .A1(n46), .A2(this_addr[1]), .ZN(n43) );
  nr03d0 U65 ( .A1(full), .A2(inc_req_n), .A3(n47), .ZN(n46) );
  inv0d0 U66 ( .I(this_addr[0]), .ZN(n47) );
endmodule


module SDRAM_FIFO_0_DW_FIFOCTL_IF_1 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [3:0] other_addr_g;
  output [3:0] word_count;
  output [2:0] this_addr;
  output [3:0] this_addr_g;
  output [3:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_3_, sync_2_, sync_1_, sync_0_, count_int_3_, empty_int, N6, N7,
         N8, N9, N10, N11, N12, N18, N19, N20, N21, N22, N23, n15, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50;

  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrn1 empty_int_reg ( .D(N18), .SD(count_int_3_), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(n15) );
  sdcrq1 count_int_reg_0_ ( .D(N6), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 count_int_reg_1_ ( .D(N7), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_2_ ( .D(N8), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_3_ ( .D(N9), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_int_3_) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N12), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N9), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N11), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N10), .SD(sync_3_), .SC(test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrq1 error_int_reg ( .D(N23), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  sdcrn1 almost_empty_int_reg ( .D(N19), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrq1 half_full_int_reg ( .D(N20), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(N21), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrq1 full_int_reg ( .D(N22), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  inv0d1 U20 ( .I(n15), .ZN(empty_int) );
  aor21d1 U25 ( .B1(empty), .B2(n20), .A(error), .Z(N23) );
  inv0d0 U26 ( .I(empty_int), .ZN(empty) );
  nr04d0 U27 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(N22) );
  aor21d1 U28 ( .B1(n21), .B2(n22), .A(n25), .Z(N21) );
  inv0d0 U29 ( .I(n26), .ZN(n22) );
  aor21d1 U30 ( .B1(n21), .B2(n24), .A(N20), .Z(N19) );
  or03d0 U31 ( .A1(n21), .A2(N20), .A3(n24), .Z(N18) );
  xn02d1 U32 ( .A1(n27), .A2(n28), .ZN(n24) );
  nd02d0 U33 ( .A1(n23), .A2(n26), .ZN(N20) );
  xn02d1 U34 ( .A1(n29), .A2(n30), .ZN(n26) );
  an02d0 U35 ( .A1(n31), .A2(n32), .Z(n30) );
  nd02d0 U36 ( .A1(n33), .A2(n34), .ZN(n29) );
  inv0d0 U37 ( .I(n25), .ZN(n23) );
  xr03d1 U38 ( .A1(sync_3_), .A2(n35), .A3(n36), .Z(n25) );
  oai221d1 U39 ( .B1(n37), .B2(n31), .C1(n37), .C2(n32), .A(n34), .ZN(n35) );
  nd02d0 U40 ( .A1(n38), .A2(n39), .ZN(n34) );
  nd02d0 U41 ( .A1(n40), .A2(n41), .ZN(n32) );
  inv0d0 U42 ( .I(n33), .ZN(n37) );
  nd02d0 U43 ( .A1(n42), .A2(N8), .ZN(n33) );
  xn02d1 U44 ( .A1(n43), .A2(n40), .ZN(n21) );
  or02d0 U45 ( .A1(n28), .A2(n27), .Z(n40) );
  xn02d1 U46 ( .A1(n44), .A2(sync_0_), .ZN(n28) );
  nd02d0 U47 ( .A1(n31), .A2(n41), .ZN(n43) );
  nd02d0 U48 ( .A1(n44), .A2(N7), .ZN(n41) );
  inv0d0 U49 ( .I(n45), .ZN(n44) );
  nd02d0 U50 ( .A1(n45), .A2(n46), .ZN(n31) );
  xn02d1 U51 ( .A1(n42), .A2(sync_1_), .ZN(n45) );
  inv0d0 U52 ( .I(n38), .ZN(n42) );
  xr02d1 U53 ( .A1(sync_3_), .A2(sync_2_), .Z(n38) );
  xr02d1 U54 ( .A1(n36), .A2(n39), .Z(N12) );
  inv0d0 U55 ( .I(N9), .ZN(n36) );
  xn02d1 U56 ( .A1(n47), .A2(count_int_3_), .ZN(N9) );
  nd02d0 U57 ( .A1(this_addr[2]), .A2(n48), .ZN(n47) );
  xr02d1 U58 ( .A1(N8), .A2(N7), .Z(N11) );
  inv0d0 U59 ( .I(n46), .ZN(N7) );
  inv0d0 U60 ( .I(n39), .ZN(N8) );
  xn02d1 U61 ( .A1(this_addr[2]), .A2(n48), .ZN(n39) );
  an12d1 U62 ( .A2(this_addr[1]), .A1(n49), .Z(n48) );
  xn02d1 U63 ( .A1(n46), .A2(N6), .ZN(N10) );
  inv0d0 U64 ( .I(n27), .ZN(N6) );
  xr02d1 U65 ( .A1(n50), .A2(this_addr[0]), .Z(n27) );
  nd02d0 U66 ( .A1(empty_int), .A2(n20), .ZN(n50) );
  xr02d1 U67 ( .A1(n49), .A2(this_addr[1]), .Z(n46) );
  nd03d0 U68 ( .A1(empty_int), .A2(n20), .A3(this_addr[0]), .ZN(n49) );
  inv0d0 U69 ( .I(inc_req_n), .ZN(n20) );
endmodule


module SDRAM_FIFO_0_DW_FIFOCTL_IF_0 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [3:0] other_addr_g;
  output [3:0] word_count;
  output [2:0] this_addr;
  output [3:0] this_addr_g;
  output [3:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_3_, sync_2_, sync_1_, sync_0_, count_int_3_, N6, N7, N8, N9, N10,
         N11, N12, N18, N19, N20, N21, N22, N23, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48;

  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrq1 full_int_reg ( .D(N22), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  sdcrq1 count_int_reg_0_ ( .D(N6), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 count_int_reg_1_ ( .D(N7), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_2_ ( .D(N8), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_3_ ( .D(N9), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_int_3_) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N9), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N12), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N11), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 half_full_int_reg ( .D(N20), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(N21), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrn1 almost_empty_int_reg ( .D(N19), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrn1 empty_int_reg ( .D(N18), .SD(count_int_3_), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(empty) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N10), .SD(sync_3_), .SC(test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrq1 error_int_reg ( .D(N23), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  aor21d1 U24 ( .B1(full), .B2(n19), .A(error), .Z(N23) );
  inv0d0 U25 ( .I(inc_req_n), .ZN(n19) );
  nr04d0 U26 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(N22) );
  aor21d1 U27 ( .B1(n20), .B2(n21), .A(n24), .Z(N21) );
  inv0d0 U28 ( .I(n25), .ZN(n21) );
  aor21d1 U29 ( .B1(n20), .B2(n23), .A(N20), .Z(N19) );
  or03d0 U30 ( .A1(n20), .A2(N20), .A3(n23), .Z(N18) );
  xn02d1 U31 ( .A1(n26), .A2(n27), .ZN(n23) );
  nd02d0 U32 ( .A1(n22), .A2(n25), .ZN(N20) );
  xn02d1 U33 ( .A1(n28), .A2(n29), .ZN(n25) );
  an12d1 U34 ( .A2(n30), .A1(n31), .Z(n29) );
  nd02d0 U35 ( .A1(n32), .A2(n33), .ZN(n28) );
  inv0d0 U36 ( .I(n24), .ZN(n22) );
  xr03d1 U37 ( .A1(sync_3_), .A2(n34), .A3(n35), .Z(n24) );
  oai221d1 U38 ( .B1(n31), .B2(n33), .C1(n31), .C2(n32), .A(n30), .ZN(n34) );
  nd02d0 U39 ( .A1(n36), .A2(N8), .ZN(n30) );
  nd02d0 U40 ( .A1(n37), .A2(n38), .ZN(n32) );
  nr02d0 U41 ( .A1(n36), .A2(N8), .ZN(n31) );
  inv0d0 U42 ( .I(n39), .ZN(N8) );
  xr02d1 U43 ( .A1(n37), .A2(n40), .Z(n20) );
  an02d0 U44 ( .A1(n38), .A2(n33), .Z(n40) );
  nd02d0 U45 ( .A1(n41), .A2(N7), .ZN(n33) );
  nd02d0 U46 ( .A1(n42), .A2(n43), .ZN(n38) );
  nd02d0 U47 ( .A1(n27), .A2(n26), .ZN(n37) );
  xn02d1 U48 ( .A1(n41), .A2(sync_0_), .ZN(n27) );
  inv0d0 U49 ( .I(n42), .ZN(n41) );
  xn02d1 U50 ( .A1(n36), .A2(sync_1_), .ZN(n42) );
  xn02d1 U51 ( .A1(sync_3_), .A2(sync_2_), .ZN(n36) );
  xr02d1 U52 ( .A1(n35), .A2(n39), .Z(N12) );
  inv0d0 U53 ( .I(N9), .ZN(n35) );
  xn02d1 U54 ( .A1(n44), .A2(count_int_3_), .ZN(N9) );
  nd02d0 U55 ( .A1(this_addr[2]), .A2(n45), .ZN(n44) );
  xn02d1 U56 ( .A1(n39), .A2(N7), .ZN(N11) );
  inv0d0 U57 ( .I(n43), .ZN(N7) );
  xn02d1 U58 ( .A1(this_addr[2]), .A2(n45), .ZN(n39) );
  an02d0 U59 ( .A1(this_addr[1]), .A2(n46), .Z(n45) );
  xr02d1 U60 ( .A1(n43), .A2(n26), .Z(N10) );
  inv0d0 U61 ( .I(N6), .ZN(n26) );
  xn02d1 U62 ( .A1(n47), .A2(n48), .ZN(N6) );
  nr02d0 U63 ( .A1(full), .A2(inc_req_n), .ZN(n48) );
  xn02d1 U64 ( .A1(n46), .A2(this_addr[1]), .ZN(n43) );
  nr03d0 U65 ( .A1(full), .A2(inc_req_n), .A3(n47), .ZN(n46) );
  inv0d0 U66 ( .I(this_addr[0]), .ZN(n47) );
endmodule


module PRGRM_CNT_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  ah01d0 U1_1_6 ( .A(A[6]), .B(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  ah01d0 U1_1_5 ( .A(A[5]), .B(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  ah01d0 U1_1_4 ( .A(A[4]), .B(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  ah01d0 U1_1_3 ( .A(A[3]), .B(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  ah01d0 U1_1_2 ( .A(A[2]), .B(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  ah01d0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry_2_), .S(SUM[1]) );
  xr02d1 U1 ( .A1(carry_7_), .A2(A[7]), .Z(SUM[7]) );
  inv0d0 U2 ( .I(A[0]), .ZN(SUM[0]) );
endmodule


module PCI_FIFO_1_DW_FIFOCTL_IF_1 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [6:0] other_addr_g;
  output [6:0] word_count;
  output [5:0] this_addr;
  output [6:0] this_addr_g;
  output [6:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_5_, sync_4_, sync_3_, sync_2_, sync_1_, sync_0_, N9, N10, N11,
         N12, N13, N14, N16, N17, N18, N19, N20, N21, N22, N30, N31, N32, N34,
         N35, count_6, other_addr_g_sync_6_, other_addr_decoded_5_,
         other_addr_decoded_4_, other_addr_decoded_3_, other_addr_decoded_2_,
         other_addr_decoded_1_, other_addr_decoded_0_, advance,
         wrd_count_p1_0_, U12_g_array_3__6_, U12_g_array_t2_2__6_,
         U12_p_array_t1_2__6_, U13_g_array_1__5_, U13_g_array_3__6_,
         U13_p_array_1__3_, U13_g_array_t1_2__6_, U13_p_array_t1_2__6_,
         U14_g_array_1__5_, U14_g_array_1__3_, U14_g_array_1__1_,
         U14_p_array_0__6_, U14_g_array_t1_0__5_, U14_g_array_t1_0__3_,
         U14_g_array_t1_0__1_, U14_g_array_t1_2__6_, U14_g_array_t2_0__5_,
         U14_g_array_t2_0__3_, U14_g_array_t2_2__6_, U14_p_array_t1_2__6_, n1,
         n30, n31, n32, n33, n34, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;

  PCI_FIFO_1_DW_inc_1 U2 ( .carry_in(advance), .a({count_6, this_addr}), 
        .carry_out(SYNOPSYS_UNCONNECTED_3), .sum({N22, N14, N13, N12, N11, N10, 
        N9}) );
  PCI_FIFO_1_DW01_sub_1 U3 ( .A({N22, N14, N13, N12, N11, N10, N9}), .B({
        other_addr_g_sync_6_, other_addr_decoded_5_, other_addr_decoded_4_, 
        other_addr_decoded_3_, other_addr_decoded_2_, other_addr_decoded_1_, 
        other_addr_decoded_0_}), .CI(1'b0), .DIFF({U14_p_array_t1_2__6_, 
        U14_g_array_t1_0__5_, U14_g_array_t2_0__5_, U14_g_array_t1_0__3_, 
        U14_g_array_t2_0__3_, U14_g_array_t1_0__1_, wrd_count_p1_0_}), .CO(
        SYNOPSYS_UNCONNECTED_4) );
  sdcrq1 sync_reg_6_ ( .D(other_addr_g[6]), .SD(sync_5_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(other_addr_g_sync_6_) );
  sdcrq1 sync_reg_5_ ( .D(other_addr_g[5]), .SD(sync_4_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_5_) );
  sdcrq1 sync_reg_4_ ( .D(other_addr_g[4]), .SD(sync_3_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_4_) );
  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrq1 count_int_reg_6_ ( .D(N22), .SD(this_addr[5]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_6) );
  sdcrq1 count_int_reg_5_ ( .D(N14), .SD(this_addr[4]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[5]) );
  sdcrq1 count_int_reg_4_ ( .D(N13), .SD(this_addr[3]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[4]) );
  sdcrq1 count_int_reg_3_ ( .D(N12), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[3]) );
  sdcrq1 count_int_reg_2_ ( .D(N11), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_1_ ( .D(N10), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_0_ ( .D(N9), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 this_addr_g_int_reg_6_ ( .D(N22), .SD(this_addr_g[5]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[6]) );
  sdcrq1 this_addr_g_int_reg_5_ ( .D(N21), .SD(this_addr_g[4]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[5]) );
  sdcrq1 this_addr_g_int_reg_4_ ( .D(N20), .SD(this_addr_g[3]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[4]) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N19), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N18), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N17), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N16), .SD(other_addr_g_sync_6_), .SC(
        test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrn1 empty_int_reg ( .D(N30), .SD(count_6), .SC(test_se), .CP(clk), .CDN(
        rst_n), .QN(empty) );
  sdcrn1 almost_empty_int_reg ( .D(N31), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrq1 half_full_int_reg ( .D(N32), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(n1), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrq1 full_int_reg ( .D(N34), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  sdcrq1 error_int_reg ( .D(N35), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  ora21d1 U6 ( .B1(U14_p_array_t1_2__6_), .B2(U14_g_array_t2_2__6_), .A(
        U14_g_array_t1_2__6_), .Z(n1) );
  nd02d0 U7 ( .A1(U14_p_array_0__6_), .A2(U14_g_array_1__5_), .ZN(
        U14_g_array_t1_2__6_) );
  nd02d0 U8 ( .A1(U14_g_array_t2_0__5_), .A2(U14_g_array_t1_0__5_), .ZN(
        U14_g_array_1__5_) );
  nr02d0 U9 ( .A1(U14_g_array_1__1_), .A2(U14_g_array_1__3_), .ZN(
        U14_g_array_t2_2__6_) );
  nd02d0 U10 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U14_g_array_1__3_) );
  inv0d0 U11 ( .I(U14_g_array_t1_0__1_), .ZN(U14_g_array_1__1_) );
  inv0d0 U12 ( .I(U13_g_array_t1_2__6_), .ZN(U13_g_array_3__6_) );
  nd02d0 U13 ( .A1(U14_p_array_0__6_), .A2(U13_g_array_1__5_), .ZN(
        U13_g_array_t1_2__6_) );
  inv0d0 U14 ( .I(U14_g_array_t1_0__5_), .ZN(U13_g_array_1__5_) );
  nr02d0 U15 ( .A1(U12_p_array_t1_2__6_), .A2(U12_g_array_t2_2__6_), .ZN(
        U12_g_array_3__6_) );
  nd02d0 U16 ( .A1(U13_p_array_1__3_), .A2(U14_g_array_1__1_), .ZN(
        U12_g_array_t2_2__6_) );
  xr02d1 U44 ( .A1(sync_0_), .A2(other_addr_decoded_1_), .Z(
        other_addr_decoded_0_) );
  xr02d1 U45 ( .A1(other_addr_decoded_2_), .A2(sync_1_), .Z(
        other_addr_decoded_1_) );
  xr02d1 U46 ( .A1(other_addr_decoded_3_), .A2(sync_2_), .Z(
        other_addr_decoded_2_) );
  xr02d1 U47 ( .A1(other_addr_decoded_4_), .A2(sync_3_), .Z(
        other_addr_decoded_3_) );
  xr02d1 U48 ( .A1(other_addr_decoded_5_), .A2(sync_4_), .Z(
        other_addr_decoded_4_) );
  xr02d1 U49 ( .A1(other_addr_g_sync_6_), .A2(sync_5_), .Z(
        other_addr_decoded_5_) );
  nr02d0 U50 ( .A1(inc_req_n), .A2(full), .ZN(advance) );
  inv0d0 U51 ( .I(n30), .ZN(U12_p_array_t1_2__6_) );
  aor21d1 U53 ( .B1(full), .B2(n31), .A(error), .Z(N35) );
  inv0d0 U54 ( .I(inc_req_n), .ZN(n31) );
  nr04d0 U55 ( .A1(n32), .A2(U14_g_array_t1_0__1_), .A3(U14_g_array_t1_0__5_), 
        .A4(U14_g_array_t2_0__5_), .ZN(N34) );
  nd03d0 U56 ( .A1(U14_p_array_t1_2__6_), .A2(n33), .A3(U13_p_array_1__3_), 
        .ZN(n32) );
  inv0d0 U57 ( .I(U13_g_array_3__6_), .ZN(N32) );
  nr02d0 U58 ( .A1(U12_g_array_3__6_), .A2(n34), .ZN(N31) );
  nd12d0 U59 ( .A1(U14_g_array_t1_0__1_), .A2(n34), .ZN(N30) );
  an03d0 U60 ( .A1(n30), .A2(n33), .A3(U13_p_array_1__3_), .Z(n34) );
  nr02d0 U61 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U13_p_array_1__3_) );
  inv0d0 U62 ( .I(wrd_count_p1_0_), .ZN(n33) );
  nr02d0 U63 ( .A1(U13_p_array_t1_2__6_), .A2(U14_g_array_t1_0__5_), .ZN(n30)
         );
  nd12d0 U64 ( .A1(U14_g_array_t2_0__5_), .A2(U14_p_array_0__6_), .ZN(
        U13_p_array_t1_2__6_) );
  inv0d0 U65 ( .I(U14_p_array_t1_2__6_), .ZN(U14_p_array_0__6_) );
  xr02d1 U66 ( .A1(N14), .A2(N22), .Z(N21) );
  xr02d1 U67 ( .A1(N14), .A2(N13), .Z(N20) );
  xr02d1 U68 ( .A1(N13), .A2(N12), .Z(N19) );
  xr02d1 U69 ( .A1(N12), .A2(N11), .Z(N18) );
  xr02d1 U70 ( .A1(N11), .A2(N10), .Z(N17) );
  xr02d1 U71 ( .A1(N10), .A2(N9), .Z(N16) );
endmodule


module PCI_FIFO_1_DW_FIFOCTL_IF_0 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si, test_so );
  input [6:0] other_addr_g;
  output [6:0] word_count;
  output [5:0] this_addr;
  output [6:0] this_addr_g;
  output [6:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error, test_so;
  wire   sync_5_, sync_4_, sync_3_, sync_2_, sync_1_, sync_0_, N9, N10, N11,
         N12, N13, N14, N16, N17, N18, N19, N20, N21, N22, N30, N31, N32, N34,
         N35, count_6, other_addr_g_sync_6_, other_addr_decoded_5_,
         other_addr_decoded_4_, other_addr_decoded_3_, other_addr_decoded_2_,
         other_addr_decoded_1_, other_addr_decoded_0_, advance,
         wrd_count_p1_0_, U12_g_array_3__6_, U12_g_array_t2_2__6_,
         U12_p_array_t1_2__6_, U13_g_array_1__5_, U13_g_array_3__6_,
         U13_p_array_1__3_, U13_g_array_t1_2__6_, U13_p_array_t1_2__6_,
         U14_g_array_1__5_, U14_g_array_1__3_, U14_g_array_1__1_,
         U14_p_array_0__6_, U14_g_array_t1_0__5_, U14_g_array_t1_0__3_,
         U14_g_array_t1_0__1_, U14_g_array_t1_2__6_, U14_g_array_t2_0__5_,
         U14_g_array_t2_0__3_, U14_g_array_t2_2__6_, U14_p_array_t1_2__6_, n1,
         n30, n31, n32, n33, n34, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;

  PCI_FIFO_1_DW_inc_0 U2 ( .carry_in(advance), .a({count_6, this_addr}), 
        .carry_out(SYNOPSYS_UNCONNECTED_3), .sum({N22, N14, N13, N12, N11, N10, 
        N9}) );
  PCI_FIFO_1_DW01_sub_0 U3 ( .A({other_addr_g_sync_6_, other_addr_decoded_5_, 
        other_addr_decoded_4_, other_addr_decoded_3_, other_addr_decoded_2_, 
        other_addr_decoded_1_, other_addr_decoded_0_}), .B({N22, N14, N13, N12, 
        N11, N10, N9}), .CI(1'b0), .DIFF({U14_p_array_t1_2__6_, 
        U14_g_array_t1_0__5_, U14_g_array_t2_0__5_, U14_g_array_t1_0__3_, 
        U14_g_array_t2_0__3_, U14_g_array_t1_0__1_, wrd_count_p1_0_}), .CO(
        SYNOPSYS_UNCONNECTED_4) );
  sdcrq1 sync_reg_6_ ( .D(other_addr_g[6]), .SD(sync_5_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(other_addr_g_sync_6_) );
  sdcrq1 sync_reg_5_ ( .D(other_addr_g[5]), .SD(sync_4_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_5_) );
  sdcrq1 sync_reg_4_ ( .D(other_addr_g[4]), .SD(sync_3_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_4_) );
  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrq1 count_int_reg_6_ ( .D(N22), .SD(this_addr[5]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_6) );
  sdcrq1 count_int_reg_5_ ( .D(N14), .SD(this_addr[4]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[5]) );
  sdcrq1 count_int_reg_4_ ( .D(N13), .SD(this_addr[3]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[4]) );
  sdcrq1 count_int_reg_3_ ( .D(N12), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[3]) );
  sdcrq1 count_int_reg_2_ ( .D(N11), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_1_ ( .D(N10), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_0_ ( .D(N9), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 this_addr_g_int_reg_6_ ( .D(N22), .SD(this_addr_g[5]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[6]) );
  sdcrq1 this_addr_g_int_reg_5_ ( .D(N21), .SD(this_addr_g[4]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[5]) );
  sdcrq1 this_addr_g_int_reg_4_ ( .D(N20), .SD(this_addr_g[3]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[4]) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N19), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N18), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N17), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N16), .SD(other_addr_g_sync_6_), .SC(
        test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrn1 empty_int_reg ( .D(N30), .SD(count_6), .SC(test_se), .CP(clk), .CDN(
        rst_n), .QN(empty) );
  sdcrq1 error_int_reg ( .D(N35), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  sdcrn1 almost_empty_int_reg ( .D(N31), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrq1 half_full_int_reg ( .D(N32), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(n1), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrq1 full_int_reg ( .D(N34), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  ora21d1 U6 ( .B1(U14_p_array_t1_2__6_), .B2(U14_g_array_t2_2__6_), .A(
        U14_g_array_t1_2__6_), .Z(n1) );
  nd02d0 U7 ( .A1(U14_p_array_0__6_), .A2(U14_g_array_1__5_), .ZN(
        U14_g_array_t1_2__6_) );
  nd02d0 U8 ( .A1(U14_g_array_t2_0__5_), .A2(U14_g_array_t1_0__5_), .ZN(
        U14_g_array_1__5_) );
  nr02d0 U9 ( .A1(U14_g_array_1__1_), .A2(U14_g_array_1__3_), .ZN(
        U14_g_array_t2_2__6_) );
  nd02d0 U10 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U14_g_array_1__3_) );
  inv0d0 U11 ( .I(U14_g_array_t1_0__1_), .ZN(U14_g_array_1__1_) );
  inv0d0 U12 ( .I(U13_g_array_t1_2__6_), .ZN(U13_g_array_3__6_) );
  nd02d0 U13 ( .A1(U14_p_array_0__6_), .A2(U13_g_array_1__5_), .ZN(
        U13_g_array_t1_2__6_) );
  inv0d0 U14 ( .I(U14_g_array_t1_0__5_), .ZN(U13_g_array_1__5_) );
  nr02d0 U15 ( .A1(U12_p_array_t1_2__6_), .A2(U12_g_array_t2_2__6_), .ZN(
        U12_g_array_3__6_) );
  nd02d0 U16 ( .A1(U13_p_array_1__3_), .A2(U14_g_array_1__1_), .ZN(
        U12_g_array_t2_2__6_) );
  xr02d1 U44 ( .A1(sync_0_), .A2(other_addr_decoded_1_), .Z(
        other_addr_decoded_0_) );
  xr02d1 U45 ( .A1(other_addr_decoded_2_), .A2(sync_1_), .Z(
        other_addr_decoded_1_) );
  xr02d1 U46 ( .A1(other_addr_decoded_3_), .A2(sync_2_), .Z(
        other_addr_decoded_2_) );
  xr02d1 U47 ( .A1(other_addr_decoded_4_), .A2(sync_3_), .Z(
        other_addr_decoded_3_) );
  xr02d1 U48 ( .A1(other_addr_decoded_5_), .A2(sync_4_), .Z(
        other_addr_decoded_4_) );
  xr02d1 U49 ( .A1(other_addr_g_sync_6_), .A2(sync_5_), .Z(
        other_addr_decoded_5_) );
  nr02d0 U50 ( .A1(inc_req_n), .A2(empty), .ZN(advance) );
  inv0d0 U51 ( .I(n30), .ZN(U12_p_array_t1_2__6_) );
  aor21d1 U53 ( .B1(empty), .B2(n31), .A(error), .Z(N35) );
  inv0d0 U54 ( .I(inc_req_n), .ZN(n31) );
  nr04d0 U55 ( .A1(n32), .A2(U14_g_array_t1_0__1_), .A3(U14_g_array_t1_0__5_), 
        .A4(U14_g_array_t2_0__5_), .ZN(N34) );
  nd03d0 U56 ( .A1(U14_p_array_t1_2__6_), .A2(n33), .A3(U13_p_array_1__3_), 
        .ZN(n32) );
  inv0d0 U57 ( .I(U13_g_array_3__6_), .ZN(N32) );
  nr02d0 U58 ( .A1(U12_g_array_3__6_), .A2(n34), .ZN(N31) );
  nd12d0 U59 ( .A1(U14_g_array_t1_0__1_), .A2(n34), .ZN(N30) );
  an03d0 U60 ( .A1(n30), .A2(n33), .A3(U13_p_array_1__3_), .Z(n34) );
  nr02d0 U61 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U13_p_array_1__3_) );
  inv0d0 U62 ( .I(wrd_count_p1_0_), .ZN(n33) );
  nr02d0 U63 ( .A1(U13_p_array_t1_2__6_), .A2(U14_g_array_t1_0__5_), .ZN(n30)
         );
  nd12d0 U64 ( .A1(U14_g_array_t2_0__5_), .A2(U14_p_array_0__6_), .ZN(
        U13_p_array_t1_2__6_) );
  inv0d0 U65 ( .I(U14_p_array_t1_2__6_), .ZN(U14_p_array_0__6_) );
  xr02d1 U66 ( .A1(N14), .A2(N22), .Z(N21) );
  xr02d1 U67 ( .A1(N14), .A2(N13), .Z(N20) );
  xr02d1 U68 ( .A1(N13), .A2(N12), .Z(N19) );
  xr02d1 U69 ( .A1(N12), .A2(N11), .Z(N18) );
  xr02d1 U70 ( .A1(N11), .A2(N10), .Z(N17) );
  xr02d1 U71 ( .A1(N10), .A2(N9), .Z(N16) );
  lanlq1 LOCKUP ( .D(this_addr_g[6]), .EN(clk), .Q(test_so) );
endmodule


module PCI_FIFO_0_DW_FIFOCTL_IF_1 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [6:0] other_addr_g;
  output [6:0] word_count;
  output [5:0] this_addr;
  output [6:0] this_addr_g;
  output [6:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_5_, sync_4_, sync_3_, sync_2_, sync_1_, sync_0_, N9, N10, N11,
         N12, N13, N14, N16, N17, N18, N19, N20, N21, N22, N30, N31, N32, N34,
         N35, count_6, other_addr_g_sync_6_, other_addr_decoded_5_,
         other_addr_decoded_4_, other_addr_decoded_3_, other_addr_decoded_2_,
         other_addr_decoded_1_, other_addr_decoded_0_, advance,
         wrd_count_p1_0_, U12_g_array_3__6_, U12_g_array_t2_2__6_,
         U12_p_array_t1_2__6_, U13_g_array_1__5_, U13_g_array_3__6_,
         U13_p_array_1__3_, U13_g_array_t1_2__6_, U13_p_array_t1_2__6_,
         U14_g_array_1__5_, U14_g_array_1__3_, U14_g_array_1__1_,
         U14_p_array_0__6_, U14_g_array_t1_0__5_, U14_g_array_t1_0__3_,
         U14_g_array_t1_0__1_, U14_g_array_t1_2__6_, U14_g_array_t2_0__5_,
         U14_g_array_t2_0__3_, U14_g_array_t2_2__6_, U14_p_array_t1_2__6_, n1,
         n30, n31, n32, n33, n34, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;

  PCI_FIFO_0_DW_inc_1 U2 ( .carry_in(advance), .a({count_6, this_addr}), 
        .carry_out(SYNOPSYS_UNCONNECTED_3), .sum({N22, N14, N13, N12, N11, N10, 
        N9}) );
  PCI_FIFO_0_DW01_sub_1 U3 ( .A({N22, N14, N13, N12, N11, N10, N9}), .B({
        other_addr_g_sync_6_, other_addr_decoded_5_, other_addr_decoded_4_, 
        other_addr_decoded_3_, other_addr_decoded_2_, other_addr_decoded_1_, 
        other_addr_decoded_0_}), .CI(1'b0), .DIFF({U14_p_array_t1_2__6_, 
        U14_g_array_t1_0__5_, U14_g_array_t2_0__5_, U14_g_array_t1_0__3_, 
        U14_g_array_t2_0__3_, U14_g_array_t1_0__1_, wrd_count_p1_0_}), .CO(
        SYNOPSYS_UNCONNECTED_4) );
  sdcrq1 sync_reg_6_ ( .D(other_addr_g[6]), .SD(sync_5_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(other_addr_g_sync_6_) );
  sdcrq1 sync_reg_5_ ( .D(other_addr_g[5]), .SD(sync_4_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_5_) );
  sdcrq1 sync_reg_4_ ( .D(other_addr_g[4]), .SD(sync_3_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_4_) );
  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrq1 count_int_reg_6_ ( .D(N22), .SD(this_addr[5]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_6) );
  sdcrq1 count_int_reg_5_ ( .D(N14), .SD(this_addr[4]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[5]) );
  sdcrq1 count_int_reg_4_ ( .D(N13), .SD(this_addr[3]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[4]) );
  sdcrq1 count_int_reg_3_ ( .D(N12), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[3]) );
  sdcrq1 count_int_reg_2_ ( .D(N11), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_1_ ( .D(N10), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_0_ ( .D(N9), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 this_addr_g_int_reg_6_ ( .D(N22), .SD(this_addr_g[5]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[6]) );
  sdcrq1 this_addr_g_int_reg_5_ ( .D(N21), .SD(this_addr_g[4]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[5]) );
  sdcrq1 this_addr_g_int_reg_4_ ( .D(N20), .SD(this_addr_g[3]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[4]) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N19), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N18), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N17), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N16), .SD(other_addr_g_sync_6_), .SC(
        test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrn1 empty_int_reg ( .D(N30), .SD(count_6), .SC(test_se), .CP(clk), .CDN(
        rst_n), .QN(empty) );
  sdcrn1 almost_empty_int_reg ( .D(N31), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrq1 half_full_int_reg ( .D(N32), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(n1), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrq1 full_int_reg ( .D(N34), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  sdcrq1 error_int_reg ( .D(N35), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  ora21d1 U6 ( .B1(U14_p_array_t1_2__6_), .B2(U14_g_array_t2_2__6_), .A(
        U14_g_array_t1_2__6_), .Z(n1) );
  nd02d0 U7 ( .A1(U14_p_array_0__6_), .A2(U14_g_array_1__5_), .ZN(
        U14_g_array_t1_2__6_) );
  nd02d0 U8 ( .A1(U14_g_array_t2_0__5_), .A2(U14_g_array_t1_0__5_), .ZN(
        U14_g_array_1__5_) );
  nr02d0 U9 ( .A1(U14_g_array_1__1_), .A2(U14_g_array_1__3_), .ZN(
        U14_g_array_t2_2__6_) );
  nd02d0 U10 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U14_g_array_1__3_) );
  inv0d0 U11 ( .I(U14_g_array_t1_0__1_), .ZN(U14_g_array_1__1_) );
  inv0d0 U12 ( .I(U13_g_array_t1_2__6_), .ZN(U13_g_array_3__6_) );
  nd02d0 U13 ( .A1(U14_p_array_0__6_), .A2(U13_g_array_1__5_), .ZN(
        U13_g_array_t1_2__6_) );
  inv0d0 U14 ( .I(U14_g_array_t1_0__5_), .ZN(U13_g_array_1__5_) );
  nr02d0 U15 ( .A1(U12_p_array_t1_2__6_), .A2(U12_g_array_t2_2__6_), .ZN(
        U12_g_array_3__6_) );
  nd02d0 U16 ( .A1(U13_p_array_1__3_), .A2(U14_g_array_1__1_), .ZN(
        U12_g_array_t2_2__6_) );
  xr02d1 U44 ( .A1(sync_0_), .A2(other_addr_decoded_1_), .Z(
        other_addr_decoded_0_) );
  xr02d1 U45 ( .A1(other_addr_decoded_2_), .A2(sync_1_), .Z(
        other_addr_decoded_1_) );
  xr02d1 U46 ( .A1(other_addr_decoded_3_), .A2(sync_2_), .Z(
        other_addr_decoded_2_) );
  xr02d1 U47 ( .A1(other_addr_decoded_4_), .A2(sync_3_), .Z(
        other_addr_decoded_3_) );
  xr02d1 U48 ( .A1(other_addr_decoded_5_), .A2(sync_4_), .Z(
        other_addr_decoded_4_) );
  xr02d1 U49 ( .A1(other_addr_g_sync_6_), .A2(sync_5_), .Z(
        other_addr_decoded_5_) );
  nr02d0 U50 ( .A1(inc_req_n), .A2(full), .ZN(advance) );
  inv0d0 U51 ( .I(n30), .ZN(U12_p_array_t1_2__6_) );
  aor21d1 U53 ( .B1(full), .B2(n31), .A(error), .Z(N35) );
  inv0d0 U54 ( .I(inc_req_n), .ZN(n31) );
  nr04d0 U55 ( .A1(n32), .A2(U14_g_array_t1_0__1_), .A3(U14_g_array_t1_0__5_), 
        .A4(U14_g_array_t2_0__5_), .ZN(N34) );
  nd03d0 U56 ( .A1(U14_p_array_t1_2__6_), .A2(n33), .A3(U13_p_array_1__3_), 
        .ZN(n32) );
  inv0d0 U57 ( .I(U13_g_array_3__6_), .ZN(N32) );
  nr02d0 U58 ( .A1(U12_g_array_3__6_), .A2(n34), .ZN(N31) );
  nd12d0 U59 ( .A1(U14_g_array_t1_0__1_), .A2(n34), .ZN(N30) );
  an03d0 U60 ( .A1(n30), .A2(n33), .A3(U13_p_array_1__3_), .Z(n34) );
  nr02d0 U61 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U13_p_array_1__3_) );
  inv0d0 U62 ( .I(wrd_count_p1_0_), .ZN(n33) );
  nr02d0 U63 ( .A1(U13_p_array_t1_2__6_), .A2(U14_g_array_t1_0__5_), .ZN(n30)
         );
  nd12d0 U64 ( .A1(U14_g_array_t2_0__5_), .A2(U14_p_array_0__6_), .ZN(
        U13_p_array_t1_2__6_) );
  inv0d0 U65 ( .I(U14_p_array_t1_2__6_), .ZN(U14_p_array_0__6_) );
  xr02d1 U66 ( .A1(N14), .A2(N22), .Z(N21) );
  xr02d1 U67 ( .A1(N14), .A2(N13), .Z(N20) );
  xr02d1 U68 ( .A1(N13), .A2(N12), .Z(N19) );
  xr02d1 U69 ( .A1(N12), .A2(N11), .Z(N18) );
  xr02d1 U70 ( .A1(N11), .A2(N10), .Z(N17) );
  xr02d1 U71 ( .A1(N10), .A2(N9), .Z(N16) );
endmodule


module PCI_FIFO_0_DW_FIFOCTL_IF_0 ( clk, rst_n, init_n, inc_req_n, 
        other_addr_g, word_count, empty, almost_empty, half_full, almost_full, 
        full, error, this_addr, this_addr_g, next_word_count, next_empty_n, 
        next_full, next_error, test, test_se, test_si );
  input [6:0] other_addr_g;
  output [6:0] word_count;
  output [5:0] this_addr;
  output [6:0] this_addr_g;
  output [6:0] next_word_count;
  input clk, rst_n, init_n, inc_req_n, test, test_se, test_si;
  output empty, almost_empty, half_full, almost_full, full, error,
         next_empty_n, next_full, next_error;
  wire   sync_5_, sync_4_, sync_3_, sync_2_, sync_1_, sync_0_, N9, N10, N11,
         N12, N13, N14, N16, N17, N18, N19, N20, N21, N22, N30, N31, N32, N34,
         N35, count_6, other_addr_g_sync_6_, other_addr_decoded_5_,
         other_addr_decoded_4_, other_addr_decoded_3_, other_addr_decoded_2_,
         other_addr_decoded_1_, other_addr_decoded_0_, advance,
         wrd_count_p1_0_, U12_g_array_3__6_, U12_g_array_t2_2__6_,
         U12_p_array_t1_2__6_, U13_g_array_1__5_, U13_g_array_3__6_,
         U13_p_array_1__3_, U13_g_array_t1_2__6_, U13_p_array_t1_2__6_,
         U14_g_array_1__5_, U14_g_array_1__3_, U14_g_array_1__1_,
         U14_p_array_0__6_, U14_g_array_t1_0__5_, U14_g_array_t1_0__3_,
         U14_g_array_t1_0__1_, U14_g_array_t1_2__6_, U14_g_array_t2_0__5_,
         U14_g_array_t2_0__3_, U14_g_array_t2_2__6_, U14_p_array_t1_2__6_, n1,
         n30, n31, n32, n33, n34, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;

  PCI_FIFO_0_DW_inc_0 U2 ( .carry_in(advance), .a({count_6, this_addr}), 
        .carry_out(SYNOPSYS_UNCONNECTED_3), .sum({N22, N14, N13, N12, N11, N10, 
        N9}) );
  PCI_FIFO_0_DW01_sub_0 U3 ( .A({other_addr_g_sync_6_, other_addr_decoded_5_, 
        other_addr_decoded_4_, other_addr_decoded_3_, other_addr_decoded_2_, 
        other_addr_decoded_1_, other_addr_decoded_0_}), .B({N22, N14, N13, N12, 
        N11, N10, N9}), .CI(1'b0), .DIFF({U14_p_array_t1_2__6_, 
        U14_g_array_t1_0__5_, U14_g_array_t2_0__5_, U14_g_array_t1_0__3_, 
        U14_g_array_t2_0__3_, U14_g_array_t1_0__1_, wrd_count_p1_0_}), .CO(
        SYNOPSYS_UNCONNECTED_4) );
  sdcrq1 sync_reg_6_ ( .D(other_addr_g[6]), .SD(sync_5_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(other_addr_g_sync_6_) );
  sdcrq1 sync_reg_5_ ( .D(other_addr_g[5]), .SD(sync_4_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_5_) );
  sdcrq1 sync_reg_4_ ( .D(other_addr_g[4]), .SD(sync_3_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_4_) );
  sdcrq1 sync_reg_3_ ( .D(other_addr_g[3]), .SD(sync_2_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_3_) );
  sdcrq1 sync_reg_2_ ( .D(other_addr_g[2]), .SD(sync_1_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_2_) );
  sdcrq1 sync_reg_1_ ( .D(other_addr_g[1]), .SD(sync_0_), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_1_) );
  sdcrq1 sync_reg_0_ ( .D(other_addr_g[0]), .SD(half_full), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(sync_0_) );
  sdcrq1 count_int_reg_6_ ( .D(N22), .SD(this_addr[5]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(count_6) );
  sdcrq1 count_int_reg_5_ ( .D(N14), .SD(this_addr[4]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[5]) );
  sdcrq1 count_int_reg_4_ ( .D(N13), .SD(this_addr[3]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[4]) );
  sdcrq1 count_int_reg_3_ ( .D(N12), .SD(this_addr[2]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[3]) );
  sdcrq1 count_int_reg_2_ ( .D(N11), .SD(this_addr[1]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[2]) );
  sdcrq1 count_int_reg_1_ ( .D(N10), .SD(this_addr[0]), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[1]) );
  sdcrq1 count_int_reg_0_ ( .D(N9), .SD(almost_full), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .Q(this_addr[0]) );
  sdcrq1 this_addr_g_int_reg_6_ ( .D(N22), .SD(this_addr_g[5]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[6]) );
  sdcrq1 this_addr_g_int_reg_5_ ( .D(N21), .SD(this_addr_g[4]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[5]) );
  sdcrq1 this_addr_g_int_reg_4_ ( .D(N20), .SD(this_addr_g[3]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[4]) );
  sdcrq1 this_addr_g_int_reg_3_ ( .D(N19), .SD(this_addr_g[2]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[3]) );
  sdcrq1 this_addr_g_int_reg_2_ ( .D(N18), .SD(this_addr_g[1]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[2]) );
  sdcrq1 this_addr_g_int_reg_1_ ( .D(N17), .SD(this_addr_g[0]), .SC(test_se), 
        .CP(clk), .CDN(rst_n), .Q(this_addr_g[1]) );
  sdcrq1 this_addr_g_int_reg_0_ ( .D(N16), .SD(other_addr_g_sync_6_), .SC(
        test_se), .CP(clk), .CDN(rst_n), .Q(this_addr_g[0]) );
  sdcrn1 empty_int_reg ( .D(N30), .SD(count_6), .SC(test_se), .CP(clk), .CDN(
        rst_n), .QN(empty) );
  sdcrq1 error_int_reg ( .D(N35), .SD(empty), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(error) );
  sdcrn1 almost_empty_int_reg ( .D(N31), .SD(test_si), .SC(test_se), .CP(clk), 
        .CDN(rst_n), .QN(almost_empty) );
  sdcrq1 half_full_int_reg ( .D(N32), .SD(full), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(half_full) );
  sdcrq1 almost_full_int_reg ( .D(n1), .SD(almost_empty), .SC(test_se), .CP(
        clk), .CDN(rst_n), .Q(almost_full) );
  sdcrq1 full_int_reg ( .D(N34), .SD(error), .SC(test_se), .CP(clk), .CDN(
        rst_n), .Q(full) );
  ora21d1 U6 ( .B1(U14_p_array_t1_2__6_), .B2(U14_g_array_t2_2__6_), .A(
        U14_g_array_t1_2__6_), .Z(n1) );
  nd02d0 U7 ( .A1(U14_p_array_0__6_), .A2(U14_g_array_1__5_), .ZN(
        U14_g_array_t1_2__6_) );
  nd02d0 U8 ( .A1(U14_g_array_t2_0__5_), .A2(U14_g_array_t1_0__5_), .ZN(
        U14_g_array_1__5_) );
  nr02d0 U9 ( .A1(U14_g_array_1__1_), .A2(U14_g_array_1__3_), .ZN(
        U14_g_array_t2_2__6_) );
  nd02d0 U10 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U14_g_array_1__3_) );
  inv0d0 U11 ( .I(U14_g_array_t1_0__1_), .ZN(U14_g_array_1__1_) );
  inv0d0 U12 ( .I(U13_g_array_t1_2__6_), .ZN(U13_g_array_3__6_) );
  nd02d0 U13 ( .A1(U14_p_array_0__6_), .A2(U13_g_array_1__5_), .ZN(
        U13_g_array_t1_2__6_) );
  inv0d0 U14 ( .I(U14_g_array_t1_0__5_), .ZN(U13_g_array_1__5_) );
  nr02d0 U15 ( .A1(U12_p_array_t1_2__6_), .A2(U12_g_array_t2_2__6_), .ZN(
        U12_g_array_3__6_) );
  nd02d0 U16 ( .A1(U13_p_array_1__3_), .A2(U14_g_array_1__1_), .ZN(
        U12_g_array_t2_2__6_) );
  xr02d1 U44 ( .A1(sync_0_), .A2(other_addr_decoded_1_), .Z(
        other_addr_decoded_0_) );
  xr02d1 U45 ( .A1(other_addr_decoded_2_), .A2(sync_1_), .Z(
        other_addr_decoded_1_) );
  xr02d1 U46 ( .A1(other_addr_decoded_3_), .A2(sync_2_), .Z(
        other_addr_decoded_2_) );
  xr02d1 U47 ( .A1(other_addr_decoded_4_), .A2(sync_3_), .Z(
        other_addr_decoded_3_) );
  xr02d1 U48 ( .A1(other_addr_decoded_5_), .A2(sync_4_), .Z(
        other_addr_decoded_4_) );
  xr02d1 U49 ( .A1(other_addr_g_sync_6_), .A2(sync_5_), .Z(
        other_addr_decoded_5_) );
  nr02d0 U50 ( .A1(inc_req_n), .A2(empty), .ZN(advance) );
  inv0d0 U51 ( .I(n30), .ZN(U12_p_array_t1_2__6_) );
  aor21d1 U53 ( .B1(empty), .B2(n31), .A(error), .Z(N35) );
  inv0d0 U54 ( .I(inc_req_n), .ZN(n31) );
  nr04d0 U55 ( .A1(n32), .A2(U14_g_array_t1_0__1_), .A3(U14_g_array_t1_0__5_), 
        .A4(U14_g_array_t2_0__5_), .ZN(N34) );
  nd03d0 U56 ( .A1(U14_p_array_t1_2__6_), .A2(n33), .A3(U13_p_array_1__3_), 
        .ZN(n32) );
  inv0d0 U57 ( .I(U13_g_array_3__6_), .ZN(N32) );
  nr02d0 U58 ( .A1(U12_g_array_3__6_), .A2(n34), .ZN(N31) );
  nd12d0 U59 ( .A1(U14_g_array_t1_0__1_), .A2(n34), .ZN(N30) );
  an03d0 U60 ( .A1(n30), .A2(n33), .A3(U13_p_array_1__3_), .Z(n34) );
  nr02d0 U61 ( .A1(U14_g_array_t2_0__3_), .A2(U14_g_array_t1_0__3_), .ZN(
        U13_p_array_1__3_) );
  inv0d0 U62 ( .I(wrd_count_p1_0_), .ZN(n33) );
  nr02d0 U63 ( .A1(U13_p_array_t1_2__6_), .A2(U14_g_array_t1_0__5_), .ZN(n30)
         );
  nd12d0 U64 ( .A1(U14_g_array_t2_0__5_), .A2(U14_p_array_0__6_), .ZN(
        U13_p_array_t1_2__6_) );
  inv0d0 U65 ( .I(U14_p_array_t1_2__6_), .ZN(U14_p_array_0__6_) );
  xr02d1 U66 ( .A1(N14), .A2(N22), .Z(N21) );
  xr02d1 U67 ( .A1(N14), .A2(N13), .Z(N20) );
  xr02d1 U68 ( .A1(N13), .A2(N12), .Z(N19) );
  xr02d1 U69 ( .A1(N12), .A2(N11), .Z(N18) );
  xr02d1 U70 ( .A1(N11), .A2(N10), .Z(N17) );
  xr02d1 U71 ( .A1(N10), .A2(N9), .Z(N16) );
endmodule


module SDRAM_FIFO_1_DW_fifoctl_s2_sf_0 ( clk_push, clk_pop, rst_n, push_req_n, 
        pop_req_n, we_n, push_empty, push_ae, push_hf, push_af, push_full, 
        push_error, pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, 
        wr_addr, rd_addr, push_word_count, pop_word_count, test, test_si1, 
        test_si2, test_se, test_so2, test_so1 );
  output [2:0] wr_addr;
  output [2:0] rd_addr;
  output [3:0] push_word_count;
  output [3:0] pop_word_count;
  input clk_push, clk_pop, rst_n, push_req_n, pop_req_n, test, test_si1,
         test_si2, test_se;
  output we_n, push_empty, push_ae, push_hf, push_af, push_full, push_error,
         pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, test_so2,
         test_so1;
  wire   rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_, wr_addr_gray_2_,
         wr_addr_gray_1_, wr_addr_gray_0_, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44;

  SDRAM_FIFO_1_DW_FIFOCTL_IF_0 U1 ( .clk(clk_push), .rst_n(rst_n), .init_n(
        1'b1), .inc_req_n(push_req_n), .other_addr_g({test_so1, 
        rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_}), .word_count({
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26}), .empty(push_empty), 
        .almost_empty(push_ae), .half_full(push_hf), .almost_full(push_af), 
        .full(push_full), .error(push_error), .this_addr(wr_addr), 
        .this_addr_g({test_so2, wr_addr_gray_2_, wr_addr_gray_1_, 
        wr_addr_gray_0_}), .next_word_count({SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30}), .next_empty_n(SYNOPSYS_UNCONNECTED_31), 
        .next_full(SYNOPSYS_UNCONNECTED_32), .next_error(
        SYNOPSYS_UNCONNECTED_33), .test(test), .test_se(test_se), .test_si(
        test_si2) );
  SDRAM_FIFO_1_DW_FIFOCTL_IF_1 U2 ( .clk(clk_pop), .rst_n(rst_n), .init_n(1'b1), .inc_req_n(pop_req_n), .other_addr_g({test_so2, wr_addr_gray_2_, 
        wr_addr_gray_1_, wr_addr_gray_0_}), .word_count({
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37}), .empty(pop_empty), 
        .almost_empty(pop_ae), .half_full(pop_hf), .almost_full(pop_af), 
        .full(pop_full), .error(pop_error), .this_addr(rd_addr), .this_addr_g(
        {test_so1, rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_}), 
        .next_word_count({SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41}), .next_empty_n(
        SYNOPSYS_UNCONNECTED_42), .next_full(SYNOPSYS_UNCONNECTED_43), 
        .next_error(SYNOPSYS_UNCONNECTED_44), .test(test), .test_se(test_se), 
        .test_si(test_si1) );
  or02d0 U6 ( .A1(push_full), .A2(push_req_n), .Z(we_n) );
endmodule


module SDRAM_FIFO_0_DW_fifoctl_s2_sf_0 ( clk_push, clk_pop, rst_n, push_req_n, 
        pop_req_n, we_n, push_empty, push_ae, push_hf, push_af, push_full, 
        push_error, pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, 
        wr_addr, rd_addr, push_word_count, pop_word_count, test, test_si1, 
        test_si2, test_se, test_so1, test_so2 );
  output [2:0] wr_addr;
  output [2:0] rd_addr;
  output [3:0] push_word_count;
  output [3:0] pop_word_count;
  input clk_push, clk_pop, rst_n, push_req_n, pop_req_n, test, test_si1,
         test_si2, test_se;
  output we_n, push_empty, push_ae, push_hf, push_af, push_full, push_error,
         pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, test_so1,
         test_so2;
  wire   rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_, wr_addr_gray_2_,
         wr_addr_gray_1_, wr_addr_gray_0_, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44;

  SDRAM_FIFO_0_DW_FIFOCTL_IF_0 U1 ( .clk(clk_push), .rst_n(rst_n), .init_n(
        1'b1), .inc_req_n(push_req_n), .other_addr_g({test_so2, 
        rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_}), .word_count({
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26}), .empty(push_empty), 
        .almost_empty(push_ae), .half_full(push_hf), .almost_full(push_af), 
        .full(push_full), .error(push_error), .this_addr(wr_addr), 
        .this_addr_g({test_so1, wr_addr_gray_2_, wr_addr_gray_1_, 
        wr_addr_gray_0_}), .next_word_count({SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30}), .next_empty_n(SYNOPSYS_UNCONNECTED_31), 
        .next_full(SYNOPSYS_UNCONNECTED_32), .next_error(
        SYNOPSYS_UNCONNECTED_33), .test(test), .test_se(test_se), .test_si(
        test_si1) );
  SDRAM_FIFO_0_DW_FIFOCTL_IF_1 U2 ( .clk(clk_pop), .rst_n(rst_n), .init_n(1'b1), .inc_req_n(pop_req_n), .other_addr_g({test_so1, wr_addr_gray_2_, 
        wr_addr_gray_1_, wr_addr_gray_0_}), .word_count({
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37}), .empty(pop_empty), 
        .almost_empty(pop_ae), .half_full(pop_hf), .almost_full(pop_af), 
        .full(pop_full), .error(pop_error), .this_addr(rd_addr), .this_addr_g(
        {test_so2, rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_}), 
        .next_word_count({SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41}), .next_empty_n(
        SYNOPSYS_UNCONNECTED_42), .next_full(SYNOPSYS_UNCONNECTED_43), 
        .next_error(SYNOPSYS_UNCONNECTED_44), .test(test), .test_se(test_se), 
        .test_si(test_si2) );
  or02d0 U6 ( .A1(push_full), .A2(push_req_n), .Z(we_n) );
endmodule


module STACK_MEM_1 ( clk, PushEnbl, PopEnbl, Stack_Full, TOS, PushDataIn, 
        PopDataOut, test_se, test_si, test_so );
  input [0:2] TOS;
  input [3:0] PushDataIn;
  output [3:0] PopDataOut;
  input clk, PushEnbl, PopEnbl, Stack_Full, test_se, test_si;
  output test_so;
  wire   N18, N19, Stack_Mem_0__3_, Stack_Mem_0__2_, Stack_Mem_0__1_,
         Stack_Mem_0__0_, Stack_Mem_1__3_, Stack_Mem_1__2_, Stack_Mem_1__1_,
         Stack_Mem_1__0_, Stack_Mem_2__3_, Stack_Mem_2__2_, Stack_Mem_2__1_,
         Stack_Mem_2__0_, Stack_Mem_3__3_, Stack_Mem_3__2_, Stack_Mem_3__1_,
         Stack_Mem_3__0_, Stack_Mem_4__3_, Stack_Mem_4__2_, Stack_Mem_4__1_,
         Stack_Mem_4__0_, Stack_Mem_5__3_, Stack_Mem_5__2_, Stack_Mem_5__1_,
         Stack_Mem_5__0_, Stack_Mem_6__3_, Stack_Mem_6__2_, Stack_Mem_6__1_,
         Stack_Mem_6__0_, Stack_Mem_7__2_, Stack_Mem_7__1_, Stack_Mem_7__0_,
         N76, N77, N78, N79, n1, n10, n15, n20, n25, n30, n35, n40, n45, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n133;

  aoi2222d1 U67 ( .A1(Stack_Mem_7__0_), .A2(n97), .B1(Stack_Mem_6__0_), .B2(
        n96), .C1(Stack_Mem_5__0_), .C2(n95), .D1(Stack_Mem_4__0_), .D2(n94), 
        .ZN(n98) );
  aoi2222d1 U68 ( .A1(Stack_Mem_3__0_), .A2(n93), .B1(Stack_Mem_2__0_), .B2(
        n92), .C1(Stack_Mem_1__0_), .C2(n91), .D1(Stack_Mem_0__0_), .D2(n90), 
        .ZN(n99) );
  aoi2222d1 U69 ( .A1(Stack_Mem_7__1_), .A2(n97), .B1(Stack_Mem_6__1_), .B2(
        n96), .C1(Stack_Mem_5__1_), .C2(n95), .D1(Stack_Mem_4__1_), .D2(n94), 
        .ZN(n88) );
  aoi2222d1 U70 ( .A1(Stack_Mem_3__1_), .A2(n93), .B1(Stack_Mem_2__1_), .B2(
        n92), .C1(Stack_Mem_1__1_), .C2(n91), .D1(Stack_Mem_0__1_), .D2(n90), 
        .ZN(n89) );
  aoi2222d1 U71 ( .A1(Stack_Mem_7__2_), .A2(n97), .B1(Stack_Mem_6__2_), .B2(
        n96), .C1(Stack_Mem_5__2_), .C2(n95), .D1(Stack_Mem_4__2_), .D2(n94), 
        .ZN(n86) );
  aoi2222d1 U72 ( .A1(Stack_Mem_3__2_), .A2(n93), .B1(Stack_Mem_2__2_), .B2(
        n92), .C1(Stack_Mem_1__2_), .C2(n91), .D1(Stack_Mem_0__2_), .D2(n90), 
        .ZN(n87) );
  aoi2222d1 U73 ( .A1(test_so), .A2(n97), .B1(Stack_Mem_6__3_), .B2(n96), .C1(
        Stack_Mem_5__3_), .C2(n95), .D1(Stack_Mem_4__3_), .D2(n94), .ZN(n84)
         );
  nr03d0 U74 ( .A1(n83), .A2(n82), .A3(n81), .ZN(n94) );
  nr03d0 U75 ( .A1(n80), .A2(n82), .A3(n81), .ZN(n95) );
  nr03d0 U76 ( .A1(n79), .A2(n82), .A3(n83), .ZN(n96) );
  nr03d0 U77 ( .A1(n79), .A2(n82), .A3(n80), .ZN(n97) );
  aoi2222d1 U78 ( .A1(Stack_Mem_3__3_), .A2(n93), .B1(Stack_Mem_2__3_), .B2(
        n92), .C1(Stack_Mem_1__3_), .C2(n91), .D1(Stack_Mem_0__3_), .D2(n90), 
        .ZN(n85) );
  nr03d0 U79 ( .A1(n81), .A2(n83), .A3(n78), .ZN(n90) );
  nr03d0 U80 ( .A1(n81), .A2(n80), .A3(n78), .ZN(n91) );
  nr03d0 U81 ( .A1(n83), .A2(n79), .A3(n78), .ZN(n92) );
  nr03d0 U82 ( .A1(n80), .A2(n79), .A3(n78), .ZN(n93) );
  aoim22d1 U83 ( .A1(N19), .A2(n77), .B1(n75), .B2(n77), .Z(n82) );
  aoim22d1 U84 ( .A1(N18), .A2(n77), .B1(n73), .B2(n77), .Z(n79) );
  aoim22d1 U85 ( .A1(n71), .A2(n77), .B1(n71), .B2(n77), .Z(n80) );
  senrq1 Stack_Mem_reg_0__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_0__2_), .ENN(
        n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__3_) );
  senrq1 Stack_Mem_reg_0__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_0__1_), .ENN(
        n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__2_) );
  senrq1 Stack_Mem_reg_0__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_0__0_), .ENN(
        n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__1_) );
  senrq1 Stack_Mem_reg_0__0_ ( .D(PushDataIn[0]), .SD(PopDataOut[3]), .ENN(n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__0_) );
  senrq1 Stack_Mem_reg_1__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_1__2_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__3_) );
  senrq1 Stack_Mem_reg_1__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_1__1_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__2_) );
  senrq1 Stack_Mem_reg_1__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_1__0_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__1_) );
  senrq1 Stack_Mem_reg_1__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_0__3_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__0_) );
  senrq1 Stack_Mem_reg_2__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_2__2_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__3_) );
  senrq1 Stack_Mem_reg_2__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_2__1_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__2_) );
  senrq1 Stack_Mem_reg_2__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_2__0_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__1_) );
  senrq1 Stack_Mem_reg_2__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_1__3_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__0_) );
  senrq1 Stack_Mem_reg_3__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_3__2_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__3_) );
  senrq1 Stack_Mem_reg_3__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_3__1_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__2_) );
  senrq1 Stack_Mem_reg_3__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_3__0_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__1_) );
  senrq1 Stack_Mem_reg_3__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_2__3_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__0_) );
  senrq1 Stack_Mem_reg_4__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_4__2_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__3_) );
  senrq1 Stack_Mem_reg_4__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_4__1_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__2_) );
  senrq1 Stack_Mem_reg_4__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_4__0_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__1_) );
  senrq1 Stack_Mem_reg_4__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_3__3_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__0_) );
  senrq1 Stack_Mem_reg_5__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_5__2_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__3_) );
  senrq1 Stack_Mem_reg_5__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_5__1_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__2_) );
  senrq1 Stack_Mem_reg_5__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_5__0_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__1_) );
  senrq1 Stack_Mem_reg_5__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_4__3_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__0_) );
  senrq1 Stack_Mem_reg_6__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_6__2_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__3_) );
  senrq1 Stack_Mem_reg_6__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_6__1_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__2_) );
  senrq1 Stack_Mem_reg_6__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_6__0_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__1_) );
  senrq1 Stack_Mem_reg_6__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_5__3_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__0_) );
  senrq1 Stack_Mem_reg_7__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_7__2_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(test_so) );
  senrq1 Stack_Mem_reg_7__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_7__1_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(Stack_Mem_7__2_) );
  senrq1 Stack_Mem_reg_7__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_7__0_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(Stack_Mem_7__1_) );
  senrq1 Stack_Mem_reg_7__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_6__3_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(Stack_Mem_7__0_) );
  senrq1 PopDataOut_reg_3_ ( .D(N76), .SD(PopDataOut[2]), .ENN(n133), .SC(
        test_se), .CP(clk), .Q(PopDataOut[3]) );
  senrq1 PopDataOut_reg_2_ ( .D(N77), .SD(PopDataOut[1]), .ENN(n133), .SC(
        test_se), .CP(clk), .Q(PopDataOut[2]) );
  senrq1 PopDataOut_reg_1_ ( .D(N78), .SD(PopDataOut[0]), .ENN(n133), .SC(
        test_se), .CP(clk), .Q(PopDataOut[1]) );
  senrq1 PopDataOut_reg_0_ ( .D(N79), .SD(test_si), .ENN(n133), .SC(test_se), 
        .CP(clk), .Q(PopDataOut[0]) );
  inv0d1 U6 ( .I(n45), .ZN(n71) );
  inv0d1 U11 ( .I(n70), .ZN(n45) );
  inv0d1 U16 ( .I(TOS[2]), .ZN(n70) );
  inv0d1 U21 ( .I(n73), .ZN(n72) );
  inv0d1 U26 ( .I(n82), .ZN(n78) );
  inv0d1 U31 ( .I(n80), .ZN(n83) );
  inv0d1 U36 ( .I(n79), .ZN(n81) );
  inv0d1 U41 ( .I(TOS[1]), .ZN(n73) );
  inv0d1 U46 ( .I(n75), .ZN(n74) );
  nd04d0 U48 ( .A1(PushEnbl), .A2(n45), .A3(n72), .A4(n74), .ZN(n1) );
  nd04d0 U49 ( .A1(PushEnbl), .A2(n45), .A3(n74), .A4(n73), .ZN(n10) );
  nd04d0 U50 ( .A1(PushEnbl), .A2(n45), .A3(n72), .A4(n75), .ZN(n15) );
  nd04d0 U51 ( .A1(PushEnbl), .A2(n45), .A3(n75), .A4(n73), .ZN(n20) );
  nd04d0 U52 ( .A1(PushEnbl), .A2(n72), .A3(n74), .A4(n71), .ZN(n25) );
  nd04d0 U53 ( .A1(PushEnbl), .A2(n74), .A3(n73), .A4(n71), .ZN(n30) );
  nd04d0 U54 ( .A1(PushEnbl), .A2(n72), .A3(n75), .A4(n71), .ZN(n35) );
  nd04d0 U55 ( .A1(PushEnbl), .A2(n75), .A3(n73), .A4(n71), .ZN(n40) );
  inv0d1 U56 ( .I(PopEnbl), .ZN(n133) );
  inv0d1 U57 ( .I(TOS[0]), .ZN(n75) );
  inv0d1 U58 ( .I(Stack_Full), .ZN(n77) );
  nd02d1 U59 ( .A1(n99), .A2(n98), .ZN(N79) );
  nd02d1 U60 ( .A1(n89), .A2(n88), .ZN(N78) );
  nd02d1 U61 ( .A1(n87), .A2(n86), .ZN(N77) );
  nd02d1 U62 ( .A1(n85), .A2(n84), .ZN(N76) );
  xr02d1 U63 ( .A1(n72), .A2(n71), .Z(N18) );
  nr02d0 U64 ( .A1(n45), .A2(n72), .ZN(n76) );
  xr02d1 U65 ( .A1(n74), .A2(n76), .Z(N19) );
endmodule


module STACK_MEM_2 ( clk, PushEnbl, PopEnbl, Stack_Full, TOS, PushDataIn, 
        PopDataOut, test_se, test_si, test_so );
  input [0:2] TOS;
  input [3:0] PushDataIn;
  output [3:0] PopDataOut;
  input clk, PushEnbl, PopEnbl, Stack_Full, test_se, test_si;
  output test_so;
  wire   N18, N19, Stack_Mem_0__3_, Stack_Mem_0__2_, Stack_Mem_0__1_,
         Stack_Mem_0__0_, Stack_Mem_1__3_, Stack_Mem_1__2_, Stack_Mem_1__1_,
         Stack_Mem_1__0_, Stack_Mem_2__3_, Stack_Mem_2__2_, Stack_Mem_2__1_,
         Stack_Mem_2__0_, Stack_Mem_3__3_, Stack_Mem_3__2_, Stack_Mem_3__1_,
         Stack_Mem_3__0_, Stack_Mem_4__3_, Stack_Mem_4__2_, Stack_Mem_4__1_,
         Stack_Mem_4__0_, Stack_Mem_5__3_, Stack_Mem_5__2_, Stack_Mem_5__1_,
         Stack_Mem_5__0_, Stack_Mem_6__3_, Stack_Mem_6__2_, Stack_Mem_6__1_,
         Stack_Mem_6__0_, Stack_Mem_7__2_, Stack_Mem_7__1_, Stack_Mem_7__0_,
         N76, N77, N78, N79, n1, n10, n15, n20, n25, n30, n35, n40, n45, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n133;

  aoi2222d1 U67 ( .A1(Stack_Mem_7__0_), .A2(n97), .B1(Stack_Mem_6__0_), .B2(
        n96), .C1(Stack_Mem_5__0_), .C2(n95), .D1(Stack_Mem_4__0_), .D2(n94), 
        .ZN(n98) );
  aoi2222d1 U68 ( .A1(Stack_Mem_3__0_), .A2(n93), .B1(Stack_Mem_2__0_), .B2(
        n92), .C1(Stack_Mem_1__0_), .C2(n91), .D1(Stack_Mem_0__0_), .D2(n90), 
        .ZN(n99) );
  aoi2222d1 U69 ( .A1(Stack_Mem_7__1_), .A2(n97), .B1(Stack_Mem_6__1_), .B2(
        n96), .C1(Stack_Mem_5__1_), .C2(n95), .D1(Stack_Mem_4__1_), .D2(n94), 
        .ZN(n88) );
  aoi2222d1 U70 ( .A1(Stack_Mem_3__1_), .A2(n93), .B1(Stack_Mem_2__1_), .B2(
        n92), .C1(Stack_Mem_1__1_), .C2(n91), .D1(Stack_Mem_0__1_), .D2(n90), 
        .ZN(n89) );
  aoi2222d1 U71 ( .A1(Stack_Mem_7__2_), .A2(n97), .B1(Stack_Mem_6__2_), .B2(
        n96), .C1(Stack_Mem_5__2_), .C2(n95), .D1(Stack_Mem_4__2_), .D2(n94), 
        .ZN(n86) );
  aoi2222d1 U72 ( .A1(Stack_Mem_3__2_), .A2(n93), .B1(Stack_Mem_2__2_), .B2(
        n92), .C1(Stack_Mem_1__2_), .C2(n91), .D1(Stack_Mem_0__2_), .D2(n90), 
        .ZN(n87) );
  aoi2222d1 U73 ( .A1(test_so), .A2(n97), .B1(Stack_Mem_6__3_), .B2(n96), .C1(
        Stack_Mem_5__3_), .C2(n95), .D1(Stack_Mem_4__3_), .D2(n94), .ZN(n84)
         );
  nr03d0 U74 ( .A1(n83), .A2(n82), .A3(n81), .ZN(n94) );
  nr03d0 U75 ( .A1(n80), .A2(n82), .A3(n81), .ZN(n95) );
  nr03d0 U76 ( .A1(n79), .A2(n82), .A3(n83), .ZN(n96) );
  nr03d0 U77 ( .A1(n79), .A2(n82), .A3(n80), .ZN(n97) );
  aoi2222d1 U78 ( .A1(Stack_Mem_3__3_), .A2(n93), .B1(Stack_Mem_2__3_), .B2(
        n92), .C1(Stack_Mem_1__3_), .C2(n91), .D1(Stack_Mem_0__3_), .D2(n90), 
        .ZN(n85) );
  nr03d0 U79 ( .A1(n81), .A2(n83), .A3(n78), .ZN(n90) );
  nr03d0 U80 ( .A1(n81), .A2(n80), .A3(n78), .ZN(n91) );
  nr03d0 U81 ( .A1(n83), .A2(n79), .A3(n78), .ZN(n92) );
  nr03d0 U82 ( .A1(n80), .A2(n79), .A3(n78), .ZN(n93) );
  aoim22d1 U83 ( .A1(N19), .A2(n77), .B1(n75), .B2(n77), .Z(n82) );
  aoim22d1 U84 ( .A1(N18), .A2(n77), .B1(n73), .B2(n77), .Z(n79) );
  aoim22d1 U85 ( .A1(n71), .A2(n77), .B1(n71), .B2(n77), .Z(n80) );
  senrq1 PopDataOut_reg_3_ ( .D(N76), .SD(PopDataOut[2]), .ENN(n133), .SC(
        test_se), .CP(clk), .Q(PopDataOut[3]) );
  senrq1 PopDataOut_reg_2_ ( .D(N77), .SD(PopDataOut[1]), .ENN(n133), .SC(
        test_se), .CP(clk), .Q(PopDataOut[2]) );
  senrq1 PopDataOut_reg_1_ ( .D(N78), .SD(PopDataOut[0]), .ENN(n133), .SC(
        test_se), .CP(clk), .Q(PopDataOut[1]) );
  senrq1 PopDataOut_reg_0_ ( .D(N79), .SD(test_si), .ENN(n133), .SC(test_se), 
        .CP(clk), .Q(PopDataOut[0]) );
  senrq1 Stack_Mem_reg_0__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_0__2_), .ENN(
        n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__3_) );
  senrq1 Stack_Mem_reg_0__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_0__1_), .ENN(
        n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__2_) );
  senrq1 Stack_Mem_reg_0__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_0__0_), .ENN(
        n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__1_) );
  senrq1 Stack_Mem_reg_0__0_ ( .D(PushDataIn[0]), .SD(PopDataOut[3]), .ENN(n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_0__0_) );
  senrq1 Stack_Mem_reg_1__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_1__2_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__3_) );
  senrq1 Stack_Mem_reg_1__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_1__1_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__2_) );
  senrq1 Stack_Mem_reg_1__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_1__0_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__1_) );
  senrq1 Stack_Mem_reg_1__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_0__3_), .ENN(
        n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_1__0_) );
  senrq1 Stack_Mem_reg_2__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_2__2_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__3_) );
  senrq1 Stack_Mem_reg_2__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_2__1_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__2_) );
  senrq1 Stack_Mem_reg_2__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_2__0_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__1_) );
  senrq1 Stack_Mem_reg_2__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_1__3_), .ENN(
        n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_2__0_) );
  senrq1 Stack_Mem_reg_3__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_3__2_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__3_) );
  senrq1 Stack_Mem_reg_3__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_3__1_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__2_) );
  senrq1 Stack_Mem_reg_3__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_3__0_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__1_) );
  senrq1 Stack_Mem_reg_3__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_2__3_), .ENN(
        n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_3__0_) );
  senrq1 Stack_Mem_reg_4__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_4__2_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__3_) );
  senrq1 Stack_Mem_reg_4__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_4__1_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__2_) );
  senrq1 Stack_Mem_reg_4__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_4__0_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__1_) );
  senrq1 Stack_Mem_reg_4__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_3__3_), .ENN(
        n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_4__0_) );
  senrq1 Stack_Mem_reg_5__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_5__2_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__3_) );
  senrq1 Stack_Mem_reg_5__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_5__1_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__2_) );
  senrq1 Stack_Mem_reg_5__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_5__0_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__1_) );
  senrq1 Stack_Mem_reg_5__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_4__3_), .ENN(
        n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_5__0_) );
  senrq1 Stack_Mem_reg_6__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_6__2_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__3_) );
  senrq1 Stack_Mem_reg_6__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_6__1_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__2_) );
  senrq1 Stack_Mem_reg_6__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_6__0_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__1_) );
  senrq1 Stack_Mem_reg_6__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_5__3_), .ENN(
        n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_6__0_) );
  senrq1 Stack_Mem_reg_7__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_7__2_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(test_so) );
  senrq1 Stack_Mem_reg_7__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_7__1_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(Stack_Mem_7__2_) );
  senrq1 Stack_Mem_reg_7__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_7__0_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(Stack_Mem_7__1_) );
  senrq1 Stack_Mem_reg_7__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_6__3_), .ENN(
        n1), .SC(test_se), .CP(clk), .Q(Stack_Mem_7__0_) );
  inv0d1 U6 ( .I(n45), .ZN(n71) );
  inv0d1 U11 ( .I(n70), .ZN(n45) );
  inv0d1 U16 ( .I(TOS[2]), .ZN(n70) );
  inv0d1 U21 ( .I(n73), .ZN(n72) );
  inv0d1 U26 ( .I(n82), .ZN(n78) );
  inv0d1 U31 ( .I(n80), .ZN(n83) );
  inv0d1 U36 ( .I(n79), .ZN(n81) );
  inv0d1 U41 ( .I(TOS[1]), .ZN(n73) );
  inv0d1 U46 ( .I(n75), .ZN(n74) );
  nd04d0 U48 ( .A1(PushEnbl), .A2(n45), .A3(n72), .A4(n74), .ZN(n1) );
  nd04d0 U49 ( .A1(PushEnbl), .A2(n45), .A3(n74), .A4(n73), .ZN(n10) );
  nd04d0 U50 ( .A1(PushEnbl), .A2(n45), .A3(n72), .A4(n75), .ZN(n15) );
  nd04d0 U51 ( .A1(PushEnbl), .A2(n45), .A3(n75), .A4(n73), .ZN(n20) );
  nd04d0 U52 ( .A1(PushEnbl), .A2(n72), .A3(n74), .A4(n71), .ZN(n25) );
  nd04d0 U53 ( .A1(PushEnbl), .A2(n74), .A3(n73), .A4(n71), .ZN(n30) );
  nd04d0 U54 ( .A1(PushEnbl), .A2(n72), .A3(n75), .A4(n71), .ZN(n35) );
  nd04d0 U55 ( .A1(PushEnbl), .A2(n75), .A3(n73), .A4(n71), .ZN(n40) );
  inv0d1 U56 ( .I(PopEnbl), .ZN(n133) );
  inv0d1 U57 ( .I(TOS[0]), .ZN(n75) );
  inv0d1 U58 ( .I(Stack_Full), .ZN(n77) );
  nd02d1 U59 ( .A1(n99), .A2(n98), .ZN(N79) );
  nd02d1 U60 ( .A1(n89), .A2(n88), .ZN(N78) );
  nd02d1 U61 ( .A1(n87), .A2(n86), .ZN(N77) );
  nd02d1 U62 ( .A1(n85), .A2(n84), .ZN(N76) );
  xr02d1 U63 ( .A1(n72), .A2(n71), .Z(N18) );
  nr02d0 U64 ( .A1(n45), .A2(n72), .ZN(n76) );
  xr02d1 U65 ( .A1(n74), .A2(n76), .Z(N19) );
endmodule


module STACK_MEM_0 ( clk, PushEnbl, PopEnbl, Stack_Full, TOS, PushDataIn, 
        PopDataOut, test_se, test_si, test_so );
  input [0:2] TOS;
  input [3:0] PushDataIn;
  output [3:0] PopDataOut;
  input clk, PushEnbl, PopEnbl, Stack_Full, test_se, test_si;
  output test_so;
  wire   N18, N19, Stack_Mem_31_, Stack_Mem_30_, Stack_Mem_29_, Stack_Mem_28_,
         Stack_Mem_27_, Stack_Mem_26_, Stack_Mem_25_, Stack_Mem_24_,
         Stack_Mem_23_, Stack_Mem_22_, Stack_Mem_21_, Stack_Mem_20_,
         Stack_Mem_19_, Stack_Mem_18_, Stack_Mem_17_, Stack_Mem_16_,
         Stack_Mem_15_, Stack_Mem_14_, Stack_Mem_13_, Stack_Mem_12_,
         Stack_Mem_11_, Stack_Mem_10_, Stack_Mem_9_, Stack_Mem_8_,
         Stack_Mem_7_, Stack_Mem_6_, Stack_Mem_5_, Stack_Mem_4_, Stack_Mem_2_,
         Stack_Mem_1_, Stack_Mem_0_, N76, N77, N78, N79, n5, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n1, n10, n15, n20, n25, n30, n35, n40,
         n45, n70, n71, n72, n73, n74, n75, n76;

  aoi2222d1 U67 ( .A1(Stack_Mem_0_), .A2(n49), .B1(Stack_Mem_4_), .B2(n50), 
        .C1(Stack_Mem_8_), .C2(n51), .D1(Stack_Mem_12_), .D2(n52), .ZN(n48) );
  aoi2222d1 U68 ( .A1(Stack_Mem_16_), .A2(n53), .B1(Stack_Mem_20_), .B2(n54), 
        .C1(Stack_Mem_24_), .C2(n55), .D1(Stack_Mem_28_), .D2(n56), .ZN(n47)
         );
  aoi2222d1 U69 ( .A1(Stack_Mem_1_), .A2(n49), .B1(Stack_Mem_5_), .B2(n50), 
        .C1(Stack_Mem_9_), .C2(n51), .D1(Stack_Mem_13_), .D2(n52), .ZN(n58) );
  aoi2222d1 U70 ( .A1(Stack_Mem_17_), .A2(n53), .B1(Stack_Mem_21_), .B2(n54), 
        .C1(Stack_Mem_25_), .C2(n55), .D1(Stack_Mem_29_), .D2(n56), .ZN(n57)
         );
  aoi2222d1 U71 ( .A1(Stack_Mem_2_), .A2(n49), .B1(Stack_Mem_6_), .B2(n50), 
        .C1(Stack_Mem_10_), .C2(n51), .D1(Stack_Mem_14_), .D2(n52), .ZN(n60)
         );
  aoi2222d1 U72 ( .A1(Stack_Mem_18_), .A2(n53), .B1(Stack_Mem_22_), .B2(n54), 
        .C1(Stack_Mem_26_), .C2(n55), .D1(Stack_Mem_30_), .D2(n56), .ZN(n59)
         );
  aoi2222d1 U73 ( .A1(test_so), .A2(n49), .B1(Stack_Mem_7_), .B2(n50), .C1(
        Stack_Mem_11_), .C2(n51), .D1(Stack_Mem_15_), .D2(n52), .ZN(n62) );
  nr03d0 U74 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n52) );
  nr03d0 U75 ( .A1(n66), .A2(n64), .A3(n65), .ZN(n51) );
  nr03d0 U76 ( .A1(n67), .A2(n64), .A3(n63), .ZN(n50) );
  nr03d0 U77 ( .A1(n67), .A2(n64), .A3(n66), .ZN(n49) );
  aoi2222d1 U78 ( .A1(Stack_Mem_19_), .A2(n53), .B1(Stack_Mem_23_), .B2(n54), 
        .C1(Stack_Mem_27_), .C2(n55), .D1(Stack_Mem_31_), .D2(n56), .ZN(n61)
         );
  nr03d0 U79 ( .A1(n65), .A2(n63), .A3(n68), .ZN(n56) );
  nr03d0 U80 ( .A1(n65), .A2(n66), .A3(n68), .ZN(n55) );
  nr03d0 U81 ( .A1(n63), .A2(n67), .A3(n68), .ZN(n54) );
  nr03d0 U82 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n53) );
  aoim22d1 U83 ( .A1(N19), .A2(n69), .B1(n75), .B2(n69), .Z(n64) );
  aoim22d1 U84 ( .A1(N18), .A2(n69), .B1(n73), .B2(n69), .Z(n67) );
  aoim22d1 U85 ( .A1(n71), .A2(n69), .B1(n71), .B2(n69), .Z(n66) );
  senrq1 PopDataOut_reg_3_ ( .D(N76), .SD(PopDataOut[2]), .ENN(n5), .SC(
        test_se), .CP(clk), .Q(PopDataOut[3]) );
  senrq1 PopDataOut_reg_2_ ( .D(N77), .SD(PopDataOut[1]), .ENN(n5), .SC(
        test_se), .CP(clk), .Q(PopDataOut[2]) );
  senrq1 PopDataOut_reg_1_ ( .D(N78), .SD(PopDataOut[0]), .ENN(n5), .SC(
        test_se), .CP(clk), .Q(PopDataOut[1]) );
  senrq1 PopDataOut_reg_0_ ( .D(N79), .SD(test_si), .ENN(n5), .SC(test_se), 
        .CP(clk), .Q(PopDataOut[0]) );
  senrq1 Stack_Mem_reg_0__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_30_), .ENN(n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_31_) );
  senrq1 Stack_Mem_reg_0__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_29_), .ENN(n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_30_) );
  senrq1 Stack_Mem_reg_0__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_28_), .ENN(n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_29_) );
  senrq1 Stack_Mem_reg_0__0_ ( .D(PushDataIn[0]), .SD(PopDataOut[3]), .ENN(n40), .SC(test_se), .CP(clk), .Q(Stack_Mem_28_) );
  senrq1 Stack_Mem_reg_1__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_26_), .ENN(n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_27_) );
  senrq1 Stack_Mem_reg_1__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_25_), .ENN(n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_26_) );
  senrq1 Stack_Mem_reg_1__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_24_), .ENN(n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_25_) );
  senrq1 Stack_Mem_reg_1__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_31_), .ENN(n20), .SC(test_se), .CP(clk), .Q(Stack_Mem_24_) );
  senrq1 Stack_Mem_reg_2__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_22_), .ENN(n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_23_) );
  senrq1 Stack_Mem_reg_2__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_21_), .ENN(n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_22_) );
  senrq1 Stack_Mem_reg_2__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_20_), .ENN(n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_21_) );
  senrq1 Stack_Mem_reg_2__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_27_), .ENN(n35), .SC(test_se), .CP(clk), .Q(Stack_Mem_20_) );
  senrq1 Stack_Mem_reg_3__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_18_), .ENN(n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_19_) );
  senrq1 Stack_Mem_reg_3__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_17_), .ENN(n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_18_) );
  senrq1 Stack_Mem_reg_3__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_16_), .ENN(n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_17_) );
  senrq1 Stack_Mem_reg_3__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_23_), .ENN(n15), .SC(test_se), .CP(clk), .Q(Stack_Mem_16_) );
  senrq1 Stack_Mem_reg_4__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_14_), .ENN(n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_15_) );
  senrq1 Stack_Mem_reg_4__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_13_), .ENN(n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_14_) );
  senrq1 Stack_Mem_reg_4__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_12_), .ENN(n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_13_) );
  senrq1 Stack_Mem_reg_4__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_19_), .ENN(n30), .SC(test_se), .CP(clk), .Q(Stack_Mem_12_) );
  senrq1 Stack_Mem_reg_5__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_10_), .ENN(n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_11_) );
  senrq1 Stack_Mem_reg_5__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_9_), .ENN(n10), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_10_) );
  senrq1 Stack_Mem_reg_5__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_8_), .ENN(n10), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_9_) );
  senrq1 Stack_Mem_reg_5__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_15_), .ENN(n10), .SC(test_se), .CP(clk), .Q(Stack_Mem_8_) );
  senrq1 Stack_Mem_reg_6__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_6_), .ENN(n25), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_7_) );
  senrq1 Stack_Mem_reg_6__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_5_), .ENN(n25), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_6_) );
  senrq1 Stack_Mem_reg_6__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_4_), .ENN(n25), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_5_) );
  senrq1 Stack_Mem_reg_6__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_11_), .ENN(n25), .SC(test_se), .CP(clk), .Q(Stack_Mem_4_) );
  senrq1 Stack_Mem_reg_7__3_ ( .D(PushDataIn[3]), .SD(Stack_Mem_2_), .ENN(n1), 
        .SC(test_se), .CP(clk), .Q(test_so) );
  senrq1 Stack_Mem_reg_7__2_ ( .D(PushDataIn[2]), .SD(Stack_Mem_1_), .ENN(n1), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_2_) );
  senrq1 Stack_Mem_reg_7__1_ ( .D(PushDataIn[1]), .SD(Stack_Mem_0_), .ENN(n1), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_1_) );
  senrq1 Stack_Mem_reg_7__0_ ( .D(PushDataIn[0]), .SD(Stack_Mem_7_), .ENN(n1), 
        .SC(test_se), .CP(clk), .Q(Stack_Mem_0_) );
  inv0d1 U6 ( .I(n45), .ZN(n71) );
  inv0d1 U11 ( .I(n70), .ZN(n45) );
  inv0d1 U16 ( .I(TOS[2]), .ZN(n70) );
  inv0d1 U21 ( .I(n73), .ZN(n72) );
  inv0d1 U26 ( .I(n64), .ZN(n68) );
  inv0d1 U31 ( .I(n66), .ZN(n63) );
  inv0d1 U36 ( .I(n67), .ZN(n65) );
  inv0d1 U41 ( .I(TOS[1]), .ZN(n73) );
  inv0d1 U46 ( .I(n75), .ZN(n74) );
  nd04d0 U48 ( .A1(PushEnbl), .A2(n45), .A3(n72), .A4(n74), .ZN(n1) );
  nd04d0 U49 ( .A1(PushEnbl), .A2(n45), .A3(n74), .A4(n73), .ZN(n10) );
  nd04d0 U50 ( .A1(PushEnbl), .A2(n45), .A3(n72), .A4(n75), .ZN(n15) );
  nd04d0 U51 ( .A1(PushEnbl), .A2(n45), .A3(n75), .A4(n73), .ZN(n20) );
  nd04d0 U52 ( .A1(PushEnbl), .A2(n72), .A3(n74), .A4(n71), .ZN(n25) );
  nd04d0 U53 ( .A1(PushEnbl), .A2(n74), .A3(n73), .A4(n71), .ZN(n30) );
  nd04d0 U54 ( .A1(PushEnbl), .A2(n72), .A3(n75), .A4(n71), .ZN(n35) );
  nd04d0 U55 ( .A1(PushEnbl), .A2(n75), .A3(n73), .A4(n71), .ZN(n40) );
  inv0d1 U56 ( .I(PopEnbl), .ZN(n5) );
  inv0d1 U57 ( .I(TOS[0]), .ZN(n75) );
  inv0d1 U58 ( .I(Stack_Full), .ZN(n69) );
  nd02d1 U59 ( .A1(n47), .A2(n48), .ZN(N79) );
  nd02d1 U60 ( .A1(n57), .A2(n58), .ZN(N78) );
  nd02d1 U61 ( .A1(n59), .A2(n60), .ZN(N77) );
  nd02d1 U62 ( .A1(n61), .A2(n62), .ZN(N76) );
  xr02d1 U63 ( .A1(n72), .A2(n71), .Z(N18) );
  nr02d0 U64 ( .A1(n45), .A2(n72), .ZN(n76) );
  xr02d1 U65 ( .A1(n74), .A2(n76), .Z(N19) );
endmodule


module STACK_FSM ( reset_n, clk, PushEnbl, PopEnbl, TOS, STACK_FULL, test_se, 
        test_si, test_so );
  output [0:2] TOS;
  input reset_n, clk, PushEnbl, PopEnbl, test_se, test_si;
  output STACK_FULL, test_so;
  wire   n41, n42, N28, N29, N43, N44, N69, n6, n8, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n29, n30,
         n31, n32, n33, n34, n35, n36, n20, n37, n38, n39, n40;
  wire   [1:0] Next_Stack;
  wire   [0:2] Next_TOS;
  wire   [1:0] Crnt_Stack;

  sdcrn1 TOS_int_reg_2_ ( .D(Next_TOS[2]), .SD(TOS[1]), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .QN(n10) );
  sdcrn1 Crnt_Stack_reg_0_ ( .D(Next_Stack[0]), .SD(test_si), .SC(test_se), 
        .CP(clk), .CDN(reset_n), .QN(n8) );
  sdcrn1 Crnt_Stack_reg_1_ ( .D(Next_Stack[1]), .SD(n15), .SC(test_se), .CP(
        clk), .CDN(reset_n), .QN(n6) );
  an02d1 U12 ( .A1(n26), .A2(PushEnbl), .Z(n11) );
  aor211d1 U23 ( .C1(n20), .C2(n11), .A(n12), .B(n13), .Z(Next_TOS[2]) );
  aor31d1 U24 ( .B1(n14), .B2(n15), .B3(PushEnbl), .A(n16), .Z(n13) );
  nr02d0 U25 ( .A1(n17), .A2(n18), .ZN(n16) );
  aoim22d1 U26 ( .A1(n20), .A2(n19), .B1(PopEnbl), .B2(n20), .Z(n17) );
  aor221d1 U27 ( .B1(n21), .B2(n22), .C1(N28), .C2(n11), .A(n12), .Z(
        Next_TOS[1]) );
  aor22d1 U28 ( .A1(TOS[1]), .A2(n23), .B1(N43), .B2(n19), .Z(n22) );
  aor221d1 U29 ( .B1(n21), .B2(n24), .C1(N29), .C2(n11), .A(n12), .Z(
        Next_TOS[0]) );
  aor22d1 U30 ( .A1(Crnt_Stack[1]), .A2(n14), .B1(n11), .B2(n25), .Z(n12) );
  aor22d1 U31 ( .A1(TOS[0]), .A2(n23), .B1(N44), .B2(n19), .Z(n24) );
  nr02d0 U32 ( .A1(n23), .A2(n27), .ZN(n19) );
  nr02d0 U33 ( .A1(n15), .A2(n29), .ZN(n26) );
  aor211d1 U34 ( .C1(Crnt_Stack[1]), .C2(n23), .A(n30), .B(n31), .Z(
        Next_Stack[1]) );
  aor31d1 U35 ( .B1(n15), .B2(n32), .B3(PopEnbl), .A(n33), .Z(n31) );
  nr03d0 U36 ( .A1(n15), .A2(n34), .A3(n38), .ZN(n33) );
  aor211d1 U37 ( .C1(PopEnbl), .C2(n15), .A(n30), .B(n35), .Z(Next_Stack[0])
         );
  aon211d1 U38 ( .C1(Crnt_Stack[0]), .C2(n25), .B(n38), .A(n36), .ZN(n35) );
  aor211d1 U39 ( .C1(n27), .C2(PopEnbl), .A(PushEnbl), .B(n15), .Z(n36) );
  nr03d0 U40 ( .A1(TOS[0]), .A2(TOS[1]), .A3(n20), .ZN(n27) );
  aor21d1 U41 ( .B1(Crnt_Stack[1]), .B2(Crnt_Stack[0]), .A(n29), .Z(n30) );
  nr03d0 U42 ( .A1(n32), .A2(Crnt_Stack[0]), .A3(n34), .ZN(N69) );
  nd03d0 U43 ( .A1(TOS[1]), .A2(TOS[0]), .A3(TOS[2]), .ZN(n34) );
  sdcrq1 STACK_FULL_reg ( .D(N69), .SD(Crnt_Stack[1]), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(STACK_FULL) );
  sdcrq1 TOS_int_reg_1_ ( .D(Next_TOS[1]), .SD(TOS[0]), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(n41) );
  sdcrq1 TOS_int_reg_0_ ( .D(Next_TOS[0]), .SD(STACK_FULL), .SC(test_se), .CP(
        clk), .CDN(reset_n), .Q(TOS[0]) );
  inv0d1 U7 ( .I(n14), .ZN(n29) );
  inv0d0 U9 ( .I(n18), .ZN(n21) );
  nd02d1 U11 ( .A1(n26), .A2(n38), .ZN(n18) );
  nd02d1 U13 ( .A1(PushEnbl), .A2(PopEnbl), .ZN(n14) );
  inv0d1 U14 ( .I(PushEnbl), .ZN(n38) );
  inv0d1 U15 ( .I(PopEnbl), .ZN(n23) );
  inv0d1 U16 ( .I(n20), .ZN(TOS[2]) );
  inv0d1 U17 ( .I(Crnt_Stack[0]), .ZN(n15) );
  inv0d1 U18 ( .I(n34), .ZN(n25) );
  inv0d1 U19 ( .I(Crnt_Stack[1]), .ZN(n32) );
  inv0d1 U20 ( .I(n42), .ZN(n20) );
  inv0d1 U21 ( .I(n10), .ZN(n42) );
  inv0d1 U22 ( .I(n37), .ZN(TOS[1]) );
  inv0d1 U44 ( .I(n41), .ZN(n37) );
  inv0d1 U45 ( .I(n8), .ZN(Crnt_Stack[0]) );
  inv0d1 U46 ( .I(n6), .ZN(Crnt_Stack[1]) );
  an02d1 U47 ( .A1(TOS[2]), .A2(TOS[1]), .Z(n39) );
  xn02d1 U48 ( .A1(TOS[1]), .A2(n20), .ZN(N28) );
  xr02d1 U49 ( .A1(TOS[0]), .A2(n39), .Z(N29) );
  xr02d1 U50 ( .A1(TOS[1]), .A2(n20), .Z(N43) );
  nr02d0 U51 ( .A1(TOS[2]), .A2(TOS[1]), .ZN(n40) );
  xr02d1 U52 ( .A1(TOS[0]), .A2(n40), .Z(N44) );
  lanlq1 LOCKUP ( .D(n20), .EN(clk), .Q(test_so) );
endmodule


module PRGRM_CNT ( reset_n, clk, Incrmnt_PC, Ld_Brnch_Addr, Ld_Rtn_Addr, 
        Imm_Addr, Return_Addr, PC, test_se, test_si );
  input [7:0] Imm_Addr;
  input [7:0] Return_Addr;
  output [7:0] PC;
  input reset_n, clk, Incrmnt_PC, Ld_Brnch_Addr, Ld_Rtn_Addr, test_se, test_si;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N32, N34, N36, N38, N40, N42, N44,
         N46, n11, n12, n1, n9, n13;

  aor222d1 U13 ( .A1(Return_Addr[7]), .A2(n11), .B1(Imm_Addr[7]), .B2(n12), 
        .C1(N13), .C2(n13), .Z(N46) );
  aor222d1 U14 ( .A1(Return_Addr[6]), .A2(n11), .B1(Imm_Addr[6]), .B2(n1), 
        .C1(N12), .C2(n13), .Z(N44) );
  aor222d1 U15 ( .A1(Return_Addr[5]), .A2(n11), .B1(Imm_Addr[5]), .B2(n12), 
        .C1(N11), .C2(n13), .Z(N42) );
  aor222d1 U16 ( .A1(Return_Addr[4]), .A2(n11), .B1(Imm_Addr[4]), .B2(n12), 
        .C1(N10), .C2(n13), .Z(N40) );
  aor222d1 U17 ( .A1(Return_Addr[3]), .A2(n11), .B1(Imm_Addr[3]), .B2(n1), 
        .C1(N9), .C2(n13), .Z(N38) );
  aor222d1 U18 ( .A1(Return_Addr[2]), .A2(n11), .B1(Imm_Addr[2]), .B2(n1), 
        .C1(N8), .C2(n13), .Z(N36) );
  aor222d1 U19 ( .A1(Return_Addr[1]), .A2(n11), .B1(Imm_Addr[1]), .B2(n1), 
        .C1(N7), .C2(n13), .Z(N34) );
  aor222d1 U20 ( .A1(Return_Addr[0]), .A2(n11), .B1(Imm_Addr[0]), .B2(n12), 
        .C1(N6), .C2(n13), .Z(N32) );
  nr02d0 U21 ( .A1(n13), .A2(Ld_Rtn_Addr), .ZN(n12) );
  an12d1 U22 ( .A2(Ld_Rtn_Addr), .A1(n13), .Z(n11) );
  PRGRM_CNT_DW01_inc_0 add_37 ( .A(PC), .SUM({N13, N12, N11, N10, N9, N8, N7, 
        N6}) );
  secrq4 PCint_reg_7_ ( .D(N46), .SD(PC[6]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[7]) );
  secrq4 PCint_reg_6_ ( .D(N44), .SD(PC[5]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[6]) );
  secrq4 PCint_reg_1_ ( .D(N34), .SD(PC[0]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[1]) );
  secrq4 PCint_reg_2_ ( .D(N36), .SD(PC[1]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[2]) );
  secrq4 PCint_reg_3_ ( .D(N38), .SD(PC[2]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[3]) );
  secrq4 PCint_reg_4_ ( .D(N40), .SD(PC[3]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[4]) );
  secrq4 PCint_reg_5_ ( .D(N42), .SD(PC[4]), .ENN(n9), .SC(test_se), .CP(clk), 
        .CDN(reset_n), .Q(PC[5]) );
  secrq4 PCint_reg_0_ ( .D(N32), .SD(test_si), .ENN(n9), .SC(test_se), .CP(clk), .CDN(reset_n), .Q(PC[0]) );
  bufbd2 U10 ( .I(Incrmnt_PC), .Z(n13) );
  nr02d0 U12 ( .A1(n13), .A2(Ld_Rtn_Addr), .ZN(n1) );
  nr03d0 U23 ( .A1(Ld_Rtn_Addr), .A2(Ld_Brnch_Addr), .A3(n13), .ZN(n9) );
endmodule


module PRGRM_DECODE ( Zro_Flag, Carry_Flag, Neg_Flag, CurrentState, 
        Crnt_Instrn, Incrmnt_PC, Ld_Brnch_Addr, Ld_Rtn_Addr );
  input [2:0] CurrentState;
  input [31:0] Crnt_Instrn;
  input Zro_Flag, Carry_Flag, Neg_Flag;
  output Incrmnt_PC, Ld_Brnch_Addr, Ld_Rtn_Addr;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27;

  an04d1 U3 ( .A1(Crnt_Instrn[18]), .A2(Crnt_Instrn[19]), .A3(Crnt_Instrn[20]), 
        .A4(Crnt_Instrn[21]), .Z(n15) );
  an03d1 U5 ( .A1(n20), .A2(n21), .A3(n25), .Z(n19) );
  an03d1 U7 ( .A1(Crnt_Instrn[17]), .A2(n20), .A3(n25), .Z(n17) );
  an03d1 U10 ( .A1(Crnt_Instrn[16]), .A2(n21), .A3(n25), .Z(n18) );
  or03d1 U11 ( .A1(Crnt_Instrn[21]), .A2(Crnt_Instrn[23]), .A3(Crnt_Instrn[22]), .Z(n26) );
  an02d1 U13 ( .A1(Crnt_Instrn[27]), .A2(n12), .Z(Ld_Rtn_Addr) );
  nr03d0 U15 ( .A1(n8), .A2(Ld_Rtn_Addr), .A3(Ld_Brnch_Addr), .ZN(Incrmnt_PC)
         );
  nr03d0 U16 ( .A1(n9), .A2(n10), .A3(n11), .ZN(Ld_Brnch_Addr) );
  nr02d0 U17 ( .A1(Crnt_Instrn[28]), .A2(Crnt_Instrn[29]), .ZN(n10) );
  aoim22d1 U18 ( .A1(Crnt_Instrn[25]), .A2(n13), .B1(Crnt_Instrn[25]), .B2(n14), .Z(n9) );
  aoi2222d1 U19 ( .A1(n15), .A2(n16), .B1(Carry_Flag), .B2(n17), .C1(Zro_Flag), 
        .C2(n18), .D1(Neg_Flag), .D2(n19), .ZN(n14) );
  nr04d0 U20 ( .A1(Crnt_Instrn[23]), .A2(Crnt_Instrn[22]), .A3(n20), .A4(n21), 
        .ZN(n16) );
  aor222d1 U21 ( .A1(n18), .A2(n22), .B1(n17), .B2(n23), .C1(n19), .C2(n24), 
        .Z(n13) );
  nr04d0 U22 ( .A1(Crnt_Instrn[19]), .A2(Crnt_Instrn[20]), .A3(Crnt_Instrn[18]), .A4(n26), .ZN(n25) );
  nr03d0 U23 ( .A1(Crnt_Instrn[31]), .A2(Crnt_Instrn[30]), .A3(n8), .ZN(n12)
         );
  nr02d0 U24 ( .A1(CurrentState[1]), .A2(CurrentState[0]), .ZN(n27) );
  inv0d1 U2 ( .I(Neg_Flag), .ZN(n24) );
  inv0d1 U4 ( .I(Carry_Flag), .ZN(n23) );
  inv0d0 U6 ( .I(Zro_Flag), .ZN(n22) );
  inv0d1 U8 ( .I(n12), .ZN(n11) );
  inv0d1 U9 ( .I(Crnt_Instrn[17]), .ZN(n21) );
  inv0d1 U12 ( .I(Crnt_Instrn[16]), .ZN(n20) );
  nd02d1 U14 ( .A1(n27), .A2(CurrentState[2]), .ZN(n8) );
endmodule


module PRGRM_FSM ( clk, reset_n, CurrentState, test_se, test_si );
  output [2:0] CurrentState;
  input clk, reset_n, test_se, test_si;
  wire   n4;
  wire   [2:0] Next_State;

  nr23d1 U6 ( .A1(CurrentState[1]), .A2(CurrentState[0]), .A3(CurrentState[2]), 
        .ZN(Next_State[2]) );
  nr02d0 U7 ( .A1(CurrentState[2]), .A2(n4), .ZN(Next_State[1]) );
  xn02d1 U8 ( .A1(CurrentState[0]), .A2(CurrentState[1]), .ZN(n4) );
  aoi21d1 U9 ( .B1(CurrentState[1]), .B2(CurrentState[2]), .A(CurrentState[0]), 
        .ZN(Next_State[0]) );
  sdcrq1 Current_State_reg_2_ ( .D(Next_State[2]), .SD(CurrentState[1]), .SC(
        test_se), .CP(clk), .CDN(reset_n), .Q(CurrentState[2]) );
  sdcrq1 Current_State_reg_0_ ( .D(Next_State[0]), .SD(test_si), .SC(test_se), 
        .CP(clk), .CDN(reset_n), .Q(CurrentState[0]) );
  sdcrq1 Current_State_reg_1_ ( .D(Next_State[1]), .SD(CurrentState[0]), .SC(
        test_se), .CP(clk), .CDN(reset_n), .Q(CurrentState[1]) );
endmodule


module ALU_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n20, n21, n22, n24, n25, n27, n28, n29, n32, n33, n34, n36, n37, n38,
         n40, n41, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55, n56,
         n57, n58;

  nd02d1 U10 ( .A1(n21), .A2(A[2]), .ZN(n24) );
  xn02d1 U11 ( .A1(n21), .A2(n22), .ZN(SUM[2]) );
  nd02d1 U14 ( .A1(A[2]), .A2(A[3]), .ZN(n27) );
  nr02d0 U15 ( .A1(n27), .A2(n20), .ZN(n28) );
  xr02d1 U17 ( .A1(n24), .A2(n25), .Z(SUM[3]) );
  nr02d0 U21 ( .A1(n29), .A2(n32), .ZN(n33) );
  xr02d1 U22 ( .A1(n29), .A2(n32), .Z(SUM[4]) );
  nr02d0 U26 ( .A1(n29), .A2(n36), .ZN(n37) );
  xn02d1 U27 ( .A1(n33), .A2(n34), .ZN(SUM[5]) );
  nd02d1 U30 ( .A1(n37), .A2(A[6]), .ZN(n40) );
  xn02d1 U31 ( .A1(n37), .A2(n38), .ZN(SUM[6]) );
  nd02d1 U34 ( .A1(A[6]), .A2(A[7]), .ZN(n43) );
  nr02d0 U35 ( .A1(n36), .A2(n43), .ZN(n44) );
  nd02d1 U36 ( .A1(n44), .A2(n28), .ZN(n45) );
  xr02d1 U38 ( .A1(n40), .A2(n41), .Z(SUM[7]) );
  xn02d1 U42 ( .A1(n46), .A2(n47), .ZN(SUM[8]) );
  nr02d0 U46 ( .A1(n45), .A2(n52), .ZN(n53) );
  xr02d1 U47 ( .A1(n49), .A2(n50), .Z(SUM[9]) );
  ah01d0 U48 ( .A(A[10]), .B(n53), .CO(n54), .S(SUM[10]) );
  ah01d0 U49 ( .A(A[11]), .B(n54), .CO(n55), .S(SUM[11]) );
  ah01d0 U50 ( .A(A[12]), .B(n55), .CO(n56), .S(SUM[12]) );
  ah01d0 U51 ( .A(A[13]), .B(n56), .CO(n57), .S(SUM[13]) );
  ah01d0 U52 ( .A(A[14]), .B(n57), .CO(n58), .S(SUM[14]) );
  xr02d1 U53 ( .A1(n58), .A2(A[15]), .Z(SUM[15]) );
  nd02d0 U56 ( .A1(A[1]), .A2(A[0]), .ZN(n20) );
  nd02d0 U57 ( .A1(A[8]), .A2(A[9]), .ZN(n52) );
  nd02d0 U58 ( .A1(n46), .A2(A[8]), .ZN(n49) );
  inv0d0 U59 ( .I(A[8]), .ZN(n47) );
  inv0d0 U60 ( .I(A[9]), .ZN(n50) );
  inv0d0 U61 ( .I(A[4]), .ZN(n32) );
  inv0d0 U62 ( .I(A[6]), .ZN(n38) );
  inv0d0 U63 ( .I(A[2]), .ZN(n22) );
  inv0d0 U64 ( .I(A[5]), .ZN(n34) );
  inv0d0 U65 ( .I(A[0]), .ZN(SUM[0]) );
  inv0d0 U66 ( .I(A[7]), .ZN(n41) );
  inv0d0 U67 ( .I(A[3]), .ZN(n25) );
  inv0d1 U68 ( .I(n28), .ZN(n29) );
  inv0d1 U69 ( .I(n20), .ZN(n21) );
  inv0d1 U70 ( .I(n45), .ZN(n46) );
  xr02d1 U71 ( .A1(A[1]), .A2(A[0]), .Z(SUM[1]) );
  nd02d0 U72 ( .A1(A[4]), .A2(A[5]), .ZN(n36) );
endmodule


module ALU_DW01_dec_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n18, n21, n25, n26, n29, n30, n33, n34, n37, n40, n41, n42, n43, n46,
         n49, n50, n51, n52, n53, n54, n55, n85;

  or02d1 U3 ( .A1(A[0]), .A2(A[1]), .Z(n18) );
  xn02d1 U4 ( .A1(A[0]), .A2(A[1]), .ZN(SUM[1]) );
  nr02d0 U8 ( .A1(n18), .A2(A[2]), .ZN(n21) );
  xn02d1 U9 ( .A1(n18), .A2(A[2]), .ZN(SUM[2]) );
  xr02d1 U17 ( .A1(n21), .A2(A[3]), .Z(SUM[3]) );
  nd02d1 U22 ( .A1(n26), .A2(n29), .ZN(n30) );
  xr02d1 U23 ( .A1(n26), .A2(A[4]), .Z(SUM[4]) );
  nr02d0 U27 ( .A1(A[5]), .A2(A[4]), .ZN(n33) );
  nd02d1 U28 ( .A1(n26), .A2(n33), .ZN(n34) );
  nr02d0 U33 ( .A1(n34), .A2(A[6]), .ZN(n37) );
  xn02d1 U34 ( .A1(n34), .A2(A[6]), .ZN(SUM[6]) );
  nr02d0 U38 ( .A1(A[7]), .A2(A[6]), .ZN(n40) );
  nd02d1 U39 ( .A1(n40), .A2(n33), .ZN(n41) );
  nr02d0 U40 ( .A1(n41), .A2(n25), .ZN(n42) );
  xr02d1 U42 ( .A1(n37), .A2(A[7]), .Z(SUM[7]) );
  nr02d0 U46 ( .A1(n43), .A2(A[8]), .ZN(n46) );
  xn02d1 U47 ( .A1(n43), .A2(A[8]), .ZN(SUM[8]) );
  nr02d0 U51 ( .A1(A[9]), .A2(A[8]), .ZN(n49) );
  nd02d1 U52 ( .A1(n42), .A2(n49), .ZN(n50) );
  xr02d1 U53 ( .A1(n46), .A2(A[9]), .Z(SUM[9]) );
  or02d1 U54 ( .A1(n50), .A2(A[10]), .Z(n51) );
  xn02d1 U55 ( .A1(n50), .A2(A[10]), .ZN(SUM[10]) );
  or02d1 U56 ( .A1(n51), .A2(A[11]), .Z(n52) );
  xn02d1 U57 ( .A1(n51), .A2(A[11]), .ZN(SUM[11]) );
  or02d1 U58 ( .A1(n52), .A2(A[12]), .Z(n53) );
  xn02d1 U59 ( .A1(n52), .A2(A[12]), .ZN(SUM[12]) );
  or02d1 U60 ( .A1(n53), .A2(A[13]), .Z(n54) );
  xn02d1 U61 ( .A1(n53), .A2(A[13]), .ZN(SUM[13]) );
  or02d1 U62 ( .A1(n54), .A2(A[14]), .Z(n55) );
  xn02d1 U63 ( .A1(n54), .A2(A[14]), .ZN(SUM[14]) );
  xn02d1 U64 ( .A1(n55), .A2(A[15]), .ZN(SUM[15]) );
  inv0d0 U67 ( .I(A[4]), .ZN(n29) );
  inv0d0 U68 ( .I(A[0]), .ZN(SUM[0]) );
  inv0d1 U69 ( .I(n25), .ZN(n26) );
  inv0d1 U70 ( .I(n42), .ZN(n43) );
  or02d1 U71 ( .A1(n85), .A2(n18), .Z(n25) );
  or02d1 U72 ( .A1(A[3]), .A2(A[2]), .Z(n85) );
  xn02d1 U73 ( .A1(n30), .A2(A[5]), .ZN(SUM[5]) );
endmodule


module ALU_DW01_add_2 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n22, n23, n27, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n67, n68, n69, n70,
         n72, n74, n76, n77, n78, n79, n80, n81, n82, n84, n85, n86, n87, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n139, n140, n141,
         n142, n143, n144, n145;

  nd02d1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(n29) );
  nd02d1 U6 ( .A1(A[1]), .A2(B[1]), .ZN(n31) );
  nr02d0 U7 ( .A1(A[1]), .A2(B[1]), .ZN(n32) );
  oai21d1 U10 ( .B1(n32), .B2(n29), .A(n31), .ZN(n33) );
  xr02d1 U12 ( .A1(n89), .A2(n29), .Z(SUM[1]) );
  nd02d1 U13 ( .A1(A[2]), .A2(B[2]), .ZN(n35) );
  nr02d0 U14 ( .A1(A[2]), .A2(B[2]), .ZN(n36) );
  oai21d1 U17 ( .B1(n34), .B2(n36), .A(n35), .ZN(n37) );
  xr02d1 U18 ( .A1(n34), .A2(n90), .Z(SUM[2]) );
  nd02d1 U19 ( .A1(A[3]), .A2(B[3]), .ZN(n38) );
  nr02d0 U20 ( .A1(A[3]), .A2(B[3]), .ZN(n39) );
  oai21d1 U23 ( .B1(n39), .B2(n35), .A(n38), .ZN(n40) );
  nr02d0 U24 ( .A1(n36), .A2(n39), .ZN(n41) );
  xn02d1 U27 ( .A1(n37), .A2(n91), .ZN(SUM[3]) );
  nr02d0 U29 ( .A1(A[4]), .A2(B[4]), .ZN(n45) );
  xn02d1 U35 ( .A1(n43), .A2(n92), .ZN(SUM[4]) );
  nr02d0 U37 ( .A1(A[5]), .A2(B[5]), .ZN(n50) );
  nd02d1 U39 ( .A1(n22), .A2(n49), .ZN(n93) );
  oai21d1 U40 ( .B1(n50), .B2(n44), .A(n49), .ZN(n51) );
  nr02d0 U41 ( .A1(n45), .A2(n50), .ZN(n52) );
  xr02d1 U43 ( .A1(n48), .A2(n93), .Z(SUM[5]) );
  nd02d1 U44 ( .A1(A[6]), .A2(B[6]), .ZN(n54) );
  nr02d0 U45 ( .A1(A[6]), .A2(B[6]), .ZN(n55) );
  nd02d1 U47 ( .A1(n23), .A2(n54), .ZN(n94) );
  oai21d1 U48 ( .B1(n53), .B2(n55), .A(n54), .ZN(n56) );
  xr02d1 U49 ( .A1(n53), .A2(n94), .Z(SUM[6]) );
  nd02d1 U50 ( .A1(A[7]), .A2(B[7]), .ZN(n57) );
  nr02d0 U51 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  oai21d1 U54 ( .B1(n58), .B2(n54), .A(n57), .ZN(n59) );
  nr02d0 U55 ( .A1(n55), .A2(n58), .ZN(n60) );
  nd02d1 U57 ( .A1(n52), .A2(n60), .ZN(n62) );
  oai21d1 U58 ( .B1(n42), .B2(n62), .A(n61), .ZN(n63) );
  xn02d1 U60 ( .A1(n56), .A2(n95), .ZN(SUM[7]) );
  nd02d1 U61 ( .A1(A[8]), .A2(B[8]), .ZN(n69) );
  nr02d0 U62 ( .A1(A[8]), .A2(B[8]), .ZN(n70) );
  xr02d1 U70 ( .A1(n64), .A2(n96), .Z(SUM[8]) );
  nd02d1 U71 ( .A1(A[9]), .A2(B[9]), .ZN(n72) );
  nd02d1 U74 ( .A1(n145), .A2(n72), .ZN(n97) );
  oai21d1 U79 ( .B1(n64), .B2(n77), .A(n76), .ZN(n78) );
  nd02d1 U81 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  nr02d0 U82 ( .A1(A[10]), .A2(B[10]), .ZN(n80) );
  nd02d1 U84 ( .A1(n27), .A2(n79), .ZN(n98) );
  oai21d1 U85 ( .B1(n76), .B2(n80), .A(n79), .ZN(n81) );
  nr02d0 U86 ( .A1(n77), .A2(n80), .ZN(n82) );
  xn02d1 U88 ( .A1(n78), .A2(n98), .ZN(SUM[10]) );
  xr02d1 U94 ( .A1(A[15]), .A2(B[15]), .Z(n99) );
  xr02d1 U95 ( .A1(n87), .A2(n99), .Z(SUM[15]) );
  ad01d2 U99 ( .A(B[12]), .B(A[12]), .CI(n84), .CO(n85), .S(SUM[12]) );
  ad01d0 U100 ( .A(B[11]), .B(A[11]), .CI(n144), .CO(n84), .S(SUM[11]) );
  or02d1 U101 ( .A1(A[0]), .A2(B[0]), .Z(n139) );
  ad01d0 U102 ( .A(B[13]), .B(A[13]), .CI(n85), .CO(n86), .S(SUM[13]) );
  nd02d0 U103 ( .A1(n86), .A2(A[14]), .ZN(n140) );
  nd02d0 U104 ( .A1(n86), .A2(B[14]), .ZN(n141) );
  xr03d1 U105 ( .A1(n86), .A2(B[14]), .A3(A[14]), .Z(SUM[14]) );
  nd02d1 U106 ( .A1(A[14]), .A2(B[14]), .ZN(n142) );
  nd03d0 U107 ( .A1(n140), .A2(n141), .A3(n142), .ZN(n87) );
  inv0d0 U108 ( .I(n42), .ZN(n43) );
  inv0d0 U109 ( .I(n63), .ZN(n64) );
  nd02d0 U110 ( .A1(n47), .A2(n44), .ZN(n92) );
  nd02d0 U111 ( .A1(n68), .A2(n145), .ZN(n77) );
  xr02d1 U112 ( .A1(n143), .A2(n97), .Z(SUM[9]) );
  ora21d1 U113 ( .B1(n64), .B2(n70), .A(n69), .Z(n143) );
  nd02d0 U114 ( .A1(n68), .A2(n69), .ZN(n96) );
  inv0d0 U115 ( .I(n50), .ZN(n22) );
  nd12d0 U116 ( .A1(n32), .A2(n31), .ZN(n89) );
  inv0d0 U117 ( .I(n44), .ZN(n46) );
  aoi21d1 U118 ( .B1(n43), .B2(n52), .A(n51), .ZN(n53) );
  inv0d1 U119 ( .I(n80), .ZN(n27) );
  aoi21d1 U120 ( .B1(n51), .B2(n60), .A(n59), .ZN(n61) );
  inv0d1 U121 ( .I(n70), .ZN(n68) );
  aoi21d1 U122 ( .B1(n33), .B2(n41), .A(n40), .ZN(n42) );
  aoi21d1 U123 ( .B1(n145), .B2(n67), .A(n74), .ZN(n76) );
  inv0d1 U124 ( .I(n72), .ZN(n74) );
  inv0d1 U125 ( .I(n69), .ZN(n67) );
  nd12d0 U126 ( .A1(n39), .A2(n38), .ZN(n91) );
  nd12d0 U127 ( .A1(n58), .A2(n57), .ZN(n95) );
  nd12d0 U128 ( .A1(n36), .A2(n35), .ZN(n90) );
  inv0d1 U129 ( .I(n55), .ZN(n23) );
  aoi21d1 U130 ( .B1(n43), .B2(n47), .A(n46), .ZN(n48) );
  inv0d1 U131 ( .I(n45), .ZN(n47) );
  nd02d1 U132 ( .A1(A[4]), .A2(B[4]), .ZN(n44) );
  aor21d1 U133 ( .B1(n63), .B2(n82), .A(n81), .Z(n144) );
  or02d1 U134 ( .A1(A[9]), .A2(B[9]), .Z(n145) );
  an02d1 U135 ( .A1(n139), .A2(n29), .Z(SUM[0]) );
  inv0d1 U136 ( .I(n33), .ZN(n34) );
  nd02d0 U137 ( .A1(A[5]), .A2(B[5]), .ZN(n49) );
endmodule


module ALU_DW01_add_3 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n19, n21, n22, n23, n26, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n65, n66,
         n67, n68, n69, n70, n72, n74, n75, n76, n77, n78, n79, n80, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n136,
         n137, n138, n139, n140;

  nr02d0 U1 ( .A1(A[0]), .A2(B[0]), .ZN(n28) );
  xn02d1 U2 ( .A1(A[0]), .A2(B[0]), .ZN(SUM[0]) );
  nd02d1 U3 ( .A1(A[1]), .A2(B[1]), .ZN(n29) );
  nr02d0 U4 ( .A1(A[1]), .A2(B[1]), .ZN(n30) );
  oai21d1 U7 ( .B1(n30), .B2(n28), .A(n29), .ZN(n31) );
  xr02d1 U9 ( .A1(n86), .A2(n28), .Z(SUM[1]) );
  nd02d1 U10 ( .A1(A[2]), .A2(B[2]), .ZN(n33) );
  nr02d0 U11 ( .A1(A[2]), .A2(B[2]), .ZN(n34) );
  oai21d1 U14 ( .B1(n32), .B2(n34), .A(n33), .ZN(n35) );
  xr02d1 U15 ( .A1(n32), .A2(n87), .Z(SUM[2]) );
  nd02d1 U16 ( .A1(A[3]), .A2(B[3]), .ZN(n36) );
  nr02d0 U17 ( .A1(A[3]), .A2(B[3]), .ZN(n37) );
  nd02d1 U19 ( .A1(n19), .A2(n36), .ZN(n88) );
  oai21d1 U20 ( .B1(n37), .B2(n33), .A(n36), .ZN(n38) );
  nr02d0 U21 ( .A1(n34), .A2(n37), .ZN(n39) );
  xn02d1 U24 ( .A1(n35), .A2(n88), .ZN(SUM[3]) );
  nd02d1 U25 ( .A1(A[4]), .A2(B[4]), .ZN(n42) );
  nr02d0 U26 ( .A1(A[4]), .A2(B[4]), .ZN(n43) );
  xn02d1 U32 ( .A1(n41), .A2(n89), .ZN(SUM[4]) );
  nr02d0 U34 ( .A1(A[5]), .A2(B[5]), .ZN(n48) );
  nd02d1 U36 ( .A1(n21), .A2(n47), .ZN(n90) );
  oai21d1 U37 ( .B1(n48), .B2(n42), .A(n47), .ZN(n49) );
  nr02d0 U38 ( .A1(n43), .A2(n48), .ZN(n50) );
  xr02d1 U40 ( .A1(n46), .A2(n90), .Z(SUM[5]) );
  nd02d1 U41 ( .A1(A[6]), .A2(B[6]), .ZN(n52) );
  nr02d0 U42 ( .A1(A[6]), .A2(B[6]), .ZN(n53) );
  nd02d1 U44 ( .A1(n22), .A2(n52), .ZN(n91) );
  oai21d1 U45 ( .B1(n51), .B2(n53), .A(n52), .ZN(n54) );
  xr02d1 U46 ( .A1(n51), .A2(n91), .Z(SUM[6]) );
  nd02d1 U47 ( .A1(A[7]), .A2(B[7]), .ZN(n55) );
  nr02d0 U48 ( .A1(A[7]), .A2(B[7]), .ZN(n56) );
  nd02d1 U50 ( .A1(n23), .A2(n55), .ZN(n92) );
  oai21d1 U51 ( .B1(n56), .B2(n52), .A(n55), .ZN(n57) );
  nr02d0 U52 ( .A1(n53), .A2(n56), .ZN(n58) );
  nd02d1 U54 ( .A1(n50), .A2(n58), .ZN(n60) );
  oai21d1 U55 ( .B1(n40), .B2(n60), .A(n59), .ZN(n61) );
  xn02d1 U57 ( .A1(n54), .A2(n92), .ZN(SUM[7]) );
  nd02d1 U58 ( .A1(A[8]), .A2(B[8]), .ZN(n67) );
  nr02d0 U59 ( .A1(A[8]), .A2(B[8]), .ZN(n68) );
  oai21d1 U66 ( .B1(n62), .B2(n68), .A(n67), .ZN(n69) );
  xr02d1 U67 ( .A1(n62), .A2(n93), .Z(SUM[8]) );
  nd02d1 U68 ( .A1(A[9]), .A2(B[9]), .ZN(n70) );
  nd02d1 U71 ( .A1(n137), .A2(n70), .ZN(n94) );
  oai21d1 U76 ( .B1(n62), .B2(n75), .A(n74), .ZN(n76) );
  xn02d1 U77 ( .A1(n69), .A2(n94), .ZN(SUM[9]) );
  nd02d1 U78 ( .A1(A[10]), .A2(B[10]), .ZN(n77) );
  nr02d0 U79 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  nd02d1 U81 ( .A1(n26), .A2(n77), .ZN(n95) );
  oai21d1 U82 ( .B1(n74), .B2(n78), .A(n77), .ZN(n79) );
  nr02d0 U83 ( .A1(n75), .A2(n78), .ZN(n80) );
  xn02d1 U85 ( .A1(n76), .A2(n95), .ZN(SUM[10]) );
  xr02d1 U91 ( .A1(A[15]), .A2(B[15]), .Z(n96) );
  xr02d1 U92 ( .A1(n85), .A2(n96), .Z(SUM[15]) );
  ad01d0 U96 ( .A(B[13]), .B(A[13]), .CI(n83), .CO(n84), .S(SUM[13]) );
  inv0d0 U97 ( .I(n40), .ZN(n41) );
  inv0d0 U98 ( .I(n61), .ZN(n62) );
  inv0d0 U99 ( .I(n31), .ZN(n32) );
  nd02d0 U100 ( .A1(n66), .A2(n67), .ZN(n93) );
  nd02d0 U101 ( .A1(n66), .A2(n137), .ZN(n75) );
  nd02d0 U102 ( .A1(n45), .A2(n42), .ZN(n89) );
  inv0d0 U103 ( .I(n48), .ZN(n21) );
  inv0d0 U104 ( .I(n37), .ZN(n19) );
  nd12d0 U105 ( .A1(n34), .A2(n33), .ZN(n87) );
  inv0d0 U106 ( .I(n42), .ZN(n44) );
  inv0d1 U107 ( .I(n68), .ZN(n66) );
  aoi21d1 U108 ( .B1(n31), .B2(n39), .A(n38), .ZN(n40) );
  aoi21d1 U109 ( .B1(n137), .B2(n65), .A(n72), .ZN(n74) );
  inv0d1 U110 ( .I(n70), .ZN(n72) );
  inv0d1 U111 ( .I(n67), .ZN(n65) );
  nd12d0 U112 ( .A1(n30), .A2(n29), .ZN(n86) );
  inv0d1 U113 ( .I(n53), .ZN(n22) );
  aoi21d1 U114 ( .B1(n41), .B2(n45), .A(n44), .ZN(n46) );
  inv0d1 U115 ( .I(n43), .ZN(n45) );
  inv0d1 U116 ( .I(n78), .ZN(n26) );
  inv0d1 U117 ( .I(n56), .ZN(n23) );
  aor21d1 U118 ( .B1(n61), .B2(n80), .A(n79), .Z(n136) );
  ad01d0 U119 ( .A(B[12]), .B(A[12]), .CI(n82), .CO(n83), .S(SUM[12]) );
  or02d1 U120 ( .A1(A[9]), .A2(B[9]), .Z(n137) );
  xr03d1 U121 ( .A1(n84), .A2(B[14]), .A3(A[14]), .Z(SUM[14]) );
  nd02d0 U122 ( .A1(n84), .A2(A[14]), .ZN(n138) );
  nd02d0 U123 ( .A1(n84), .A2(B[14]), .ZN(n139) );
  nd02d0 U124 ( .A1(A[14]), .A2(B[14]), .ZN(n140) );
  nd03d0 U125 ( .A1(n138), .A2(n139), .A3(n140), .ZN(n85) );
  aoi21d1 U126 ( .B1(n41), .B2(n50), .A(n49), .ZN(n51) );
  aoi21d1 U127 ( .B1(n49), .B2(n58), .A(n57), .ZN(n59) );
  nd02d0 U128 ( .A1(A[5]), .A2(B[5]), .ZN(n47) );
  ad01d2 U129 ( .A(B[11]), .B(A[11]), .CI(n136), .CO(n82), .S(SUM[11]) );
endmodule


module ALU_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n36, n38, n40, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n83, n84, n85,
         n86, n88, n90, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n158, n159, n160;

  nd02d1 U22 ( .A1(n18), .A2(A[1]), .ZN(n47) );
  nr02d0 U23 ( .A1(n18), .A2(A[1]), .ZN(n48) );
  oai21d1 U26 ( .B1(n48), .B2(n45), .A(n47), .ZN(n49) );
  xr02d1 U28 ( .A1(n107), .A2(n45), .Z(DIFF[1]) );
  nd02d1 U29 ( .A1(n19), .A2(A[2]), .ZN(n51) );
  nr02d0 U30 ( .A1(n19), .A2(A[2]), .ZN(n52) );
  oai21d1 U33 ( .B1(n50), .B2(n52), .A(n51), .ZN(n53) );
  xr02d1 U34 ( .A1(n50), .A2(n108), .Z(DIFF[2]) );
  nd02d1 U35 ( .A1(n20), .A2(A[3]), .ZN(n54) );
  nr02d0 U36 ( .A1(n20), .A2(A[3]), .ZN(n55) );
  nd02d1 U38 ( .A1(n36), .A2(n54), .ZN(n109) );
  oai21d1 U39 ( .B1(n55), .B2(n51), .A(n54), .ZN(n56) );
  nr02d0 U40 ( .A1(n52), .A2(n55), .ZN(n57) );
  xn02d1 U43 ( .A1(n53), .A2(n109), .ZN(DIFF[3]) );
  nr02d0 U45 ( .A1(A[4]), .A2(n21), .ZN(n61) );
  nd02d1 U47 ( .A1(n63), .A2(n60), .ZN(n110) );
  xn02d1 U51 ( .A1(n59), .A2(n110), .ZN(DIFF[4]) );
  nr02d0 U53 ( .A1(A[5]), .A2(n22), .ZN(n66) );
  nd02d1 U55 ( .A1(n38), .A2(n65), .ZN(n111) );
  oai21d1 U56 ( .B1(n66), .B2(n60), .A(n65), .ZN(n67) );
  nr02d0 U57 ( .A1(n61), .A2(n66), .ZN(n68) );
  xr02d1 U59 ( .A1(n64), .A2(n111), .Z(DIFF[5]) );
  nd02d1 U60 ( .A1(A[6]), .A2(n23), .ZN(n70) );
  nr02d0 U61 ( .A1(A[6]), .A2(n23), .ZN(n71) );
  oai21d1 U64 ( .B1(n69), .B2(n71), .A(n70), .ZN(n72) );
  xr02d1 U65 ( .A1(n69), .A2(n112), .Z(DIFF[6]) );
  nd02d1 U66 ( .A1(A[7]), .A2(n24), .ZN(n73) );
  nr02d0 U67 ( .A1(A[7]), .A2(n24), .ZN(n74) );
  nd02d1 U69 ( .A1(n40), .A2(n73), .ZN(n113) );
  oai21d1 U70 ( .B1(n74), .B2(n70), .A(n73), .ZN(n75) );
  nr02d0 U71 ( .A1(n71), .A2(n74), .ZN(n76) );
  nd02d1 U73 ( .A1(n68), .A2(n76), .ZN(n78) );
  oai21d1 U74 ( .B1(n58), .B2(n78), .A(n77), .ZN(n79) );
  xn02d1 U76 ( .A1(n72), .A2(n113), .ZN(DIFF[7]) );
  nr02d0 U78 ( .A1(A[8]), .A2(n25), .ZN(n86) );
  xr02d1 U86 ( .A1(n80), .A2(n114), .Z(DIFF[8]) );
  nd02d1 U90 ( .A1(n160), .A2(n88), .ZN(n115) );
  oai21d1 U95 ( .B1(n80), .B2(n93), .A(n92), .ZN(n94) );
  nd02d1 U97 ( .A1(A[10]), .A2(n27), .ZN(n95) );
  nr02d0 U98 ( .A1(A[10]), .A2(n27), .ZN(n96) );
  oai21d1 U101 ( .B1(n92), .B2(n96), .A(n95), .ZN(n97) );
  nr02d0 U102 ( .A1(n93), .A2(n96), .ZN(n98) );
  xn02d1 U104 ( .A1(n94), .A2(n116), .ZN(DIFF[10]) );
  nd02d1 U105 ( .A1(n28), .A2(A[11]), .ZN(n100) );
  nr02d0 U106 ( .A1(n28), .A2(A[11]), .ZN(n101) );
  oai21d1 U109 ( .B1(n99), .B2(n101), .A(n100), .ZN(n102) );
  xr02d1 U110 ( .A1(n99), .A2(n117), .Z(DIFF[11]) );
  xr02d1 U115 ( .A1(n105), .A2(n118), .Z(DIFF[15]) );
  ad01d1 U119 ( .A(A[13]), .B(n30), .CI(n103), .CO(n104), .S(DIFF[13]) );
  or02d1 U120 ( .A1(A[0]), .A2(n17), .Z(n158) );
  ad01d2 U121 ( .A(A[12]), .B(n29), .CI(n102), .CO(n103), .S(DIFF[12]) );
  nd02d0 U122 ( .A1(A[8]), .A2(n25), .ZN(n85) );
  nd02d1 U123 ( .A1(A[4]), .A2(n21), .ZN(n60) );
  nd02d1 U124 ( .A1(A[0]), .A2(n17), .ZN(n45) );
  inv0d1 U125 ( .I(B[0]), .ZN(n17) );
  ad01d0 U126 ( .A(A[14]), .B(n31), .CI(n104), .CO(n105), .S(DIFF[14]) );
  inv0d0 U127 ( .I(n58), .ZN(n59) );
  inv0d0 U128 ( .I(n79), .ZN(n80) );
  inv0d0 U129 ( .I(n49), .ZN(n50) );
  nd02d0 U130 ( .A1(n84), .A2(n160), .ZN(n93) );
  nd02d0 U131 ( .A1(n84), .A2(n85), .ZN(n114) );
  xr02d1 U132 ( .A1(n159), .A2(n115), .Z(DIFF[9]) );
  ora21d1 U133 ( .B1(n80), .B2(n86), .A(n85), .Z(n159) );
  inv0d0 U134 ( .I(n74), .ZN(n40) );
  nd12d0 U135 ( .A1(n71), .A2(n70), .ZN(n112) );
  inv0d0 U136 ( .I(n66), .ZN(n38) );
  nd12d0 U137 ( .A1(n52), .A2(n51), .ZN(n108) );
  inv0d0 U138 ( .I(n55), .ZN(n36) );
  inv0d0 U139 ( .I(n60), .ZN(n62) );
  nd02d0 U140 ( .A1(A[9]), .A2(n26), .ZN(n88) );
  inv0d0 U141 ( .I(B[6]), .ZN(n23) );
  inv0d0 U142 ( .I(B[2]), .ZN(n19) );
  inv0d0 U143 ( .I(B[7]), .ZN(n24) );
  aoi21d1 U144 ( .B1(n59), .B2(n68), .A(n67), .ZN(n69) );
  aoi21d1 U145 ( .B1(n67), .B2(n76), .A(n75), .ZN(n77) );
  inv0d1 U146 ( .I(n86), .ZN(n84) );
  aoi21d1 U147 ( .B1(n49), .B2(n57), .A(n56), .ZN(n58) );
  aoi21d1 U148 ( .B1(n79), .B2(n98), .A(n97), .ZN(n99) );
  aoi21d1 U149 ( .B1(n160), .B2(n83), .A(n90), .ZN(n92) );
  inv0d1 U150 ( .I(n88), .ZN(n90) );
  inv0d1 U151 ( .I(n85), .ZN(n83) );
  nd12d0 U152 ( .A1(n96), .A2(n95), .ZN(n116) );
  aoi21d1 U153 ( .B1(n59), .B2(n63), .A(n62), .ZN(n64) );
  inv0d1 U154 ( .I(n61), .ZN(n63) );
  nd12d0 U155 ( .A1(n48), .A2(n47), .ZN(n107) );
  or02d1 U156 ( .A1(A[9]), .A2(n26), .Z(n160) );
  nd12d0 U157 ( .A1(n101), .A2(n100), .ZN(n117) );
  an02d1 U158 ( .A1(n158), .A2(n45), .Z(DIFF[0]) );
  inv0d1 U159 ( .I(B[13]), .ZN(n30) );
  inv0d1 U160 ( .I(B[14]), .ZN(n31) );
  inv0d1 U161 ( .I(B[4]), .ZN(n21) );
  inv0d1 U162 ( .I(B[12]), .ZN(n29) );
  inv0d1 U163 ( .I(B[11]), .ZN(n28) );
  inv0d1 U164 ( .I(B[1]), .ZN(n18) );
  inv0d1 U165 ( .I(B[3]), .ZN(n20) );
  inv0d1 U166 ( .I(B[9]), .ZN(n26) );
  inv0d1 U167 ( .I(B[8]), .ZN(n25) );
  inv0d1 U168 ( .I(B[10]), .ZN(n27) );
  inv0d1 U169 ( .I(B[5]), .ZN(n22) );
  xn02d1 U170 ( .A1(B[15]), .A2(A[15]), .ZN(n118) );
  nd02d0 U171 ( .A1(A[5]), .A2(n22), .ZN(n65) );
endmodule


module ALU_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n35, n37, n39, n44, n45, n46, n47, n48, n49, n50, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n82, n83, n84, n85,
         n86, n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n155, n156, n157, n158, n159, n160;

  nr02d0 U17 ( .A1(A[0]), .A2(n17), .ZN(n44) );
  xn02d1 U18 ( .A1(A[0]), .A2(n17), .ZN(DIFF[0]) );
  nd02d1 U19 ( .A1(n18), .A2(A[1]), .ZN(n45) );
  nr02d0 U20 ( .A1(n18), .A2(A[1]), .ZN(n46) );
  oai21d1 U23 ( .B1(n46), .B2(n44), .A(n45), .ZN(n47) );
  xr02d1 U25 ( .A1(n104), .A2(n44), .Z(DIFF[1]) );
  nd02d1 U26 ( .A1(n19), .A2(A[2]), .ZN(n49) );
  nr02d0 U27 ( .A1(n19), .A2(A[2]), .ZN(n50) );
  xr02d1 U31 ( .A1(n48), .A2(n105), .Z(DIFF[2]) );
  nd02d1 U32 ( .A1(n20), .A2(A[3]), .ZN(n52) );
  nr02d0 U33 ( .A1(n20), .A2(A[3]), .ZN(n53) );
  nd02d1 U35 ( .A1(n35), .A2(n52), .ZN(n106) );
  oai21d1 U36 ( .B1(n53), .B2(n49), .A(n52), .ZN(n54) );
  nr02d0 U37 ( .A1(n50), .A2(n53), .ZN(n55) );
  nr02d0 U42 ( .A1(A[4]), .A2(n21), .ZN(n59) );
  nd02d1 U44 ( .A1(n61), .A2(n58), .ZN(n107) );
  xn02d1 U48 ( .A1(n57), .A2(n107), .ZN(DIFF[4]) );
  nr02d0 U50 ( .A1(A[5]), .A2(n22), .ZN(n64) );
  nd02d1 U52 ( .A1(n37), .A2(n63), .ZN(n108) );
  oai21d1 U53 ( .B1(n64), .B2(n58), .A(n63), .ZN(n65) );
  nr02d0 U54 ( .A1(n59), .A2(n64), .ZN(n66) );
  nd02d1 U57 ( .A1(A[6]), .A2(n23), .ZN(n68) );
  nr02d0 U58 ( .A1(A[6]), .A2(n23), .ZN(n69) );
  oai21d1 U61 ( .B1(n67), .B2(n69), .A(n68), .ZN(n70) );
  xr02d1 U62 ( .A1(n67), .A2(n109), .Z(DIFF[6]) );
  nd02d1 U63 ( .A1(A[7]), .A2(n24), .ZN(n71) );
  nr02d0 U64 ( .A1(A[7]), .A2(n24), .ZN(n72) );
  nd02d1 U66 ( .A1(n39), .A2(n71), .ZN(n110) );
  oai21d1 U67 ( .B1(n72), .B2(n68), .A(n71), .ZN(n73) );
  nr02d0 U68 ( .A1(n69), .A2(n72), .ZN(n74) );
  nd02d1 U70 ( .A1(n66), .A2(n74), .ZN(n76) );
  oai21d1 U71 ( .B1(n56), .B2(n76), .A(n75), .ZN(n77) );
  xn02d1 U73 ( .A1(n70), .A2(n110), .ZN(DIFF[7]) );
  nr02d0 U75 ( .A1(A[8]), .A2(n25), .ZN(n84) );
  oai21d1 U82 ( .B1(n78), .B2(n84), .A(n83), .ZN(n85) );
  xr02d1 U83 ( .A1(n78), .A2(n111), .Z(DIFF[8]) );
  oai21d1 U92 ( .B1(n78), .B2(n91), .A(n90), .ZN(n92) );
  xn02d1 U93 ( .A1(n85), .A2(n112), .ZN(DIFF[9]) );
  nd02d1 U94 ( .A1(A[10]), .A2(n27), .ZN(n93) );
  nr02d0 U95 ( .A1(A[10]), .A2(n27), .ZN(n94) );
  oai21d1 U98 ( .B1(n90), .B2(n94), .A(n93), .ZN(n95) );
  nr02d0 U99 ( .A1(n91), .A2(n94), .ZN(n96) );
  xn02d1 U101 ( .A1(n92), .A2(n113), .ZN(DIFF[10]) );
  nd02d1 U102 ( .A1(n28), .A2(A[11]), .ZN(n98) );
  nr02d0 U103 ( .A1(n28), .A2(A[11]), .ZN(n99) );
  oai21d1 U106 ( .B1(n97), .B2(n99), .A(n98), .ZN(n100) );
  xr02d1 U107 ( .A1(n97), .A2(n114), .Z(DIFF[11]) );
  xr02d1 U112 ( .A1(n103), .A2(n115), .Z(DIFF[15]) );
  ad01d2 U116 ( .A(A[12]), .B(n29), .CI(n100), .CO(n101), .S(DIFF[12]) );
  nd02d1 U117 ( .A1(n102), .A2(A[14]), .ZN(n155) );
  ad01d0 U118 ( .A(A[13]), .B(n30), .CI(n101), .CO(n102), .S(DIFF[13]) );
  inv0d1 U119 ( .I(B[14]), .ZN(n31) );
  xr03d1 U120 ( .A1(n102), .A2(n31), .A3(A[14]), .Z(DIFF[14]) );
  nd02d1 U121 ( .A1(n102), .A2(n31), .ZN(n156) );
  nd02d0 U122 ( .A1(A[14]), .A2(n31), .ZN(n157) );
  nd03d0 U123 ( .A1(n155), .A2(n156), .A3(n157), .ZN(n103) );
  nd02d1 U124 ( .A1(A[8]), .A2(n25), .ZN(n83) );
  inv0d1 U125 ( .I(B[0]), .ZN(n17) );
  inv0d0 U126 ( .I(n56), .ZN(n57) );
  inv0d0 U127 ( .I(n77), .ZN(n78) );
  inv0d0 U128 ( .I(n47), .ZN(n48) );
  nd02d0 U129 ( .A1(n82), .A2(n160), .ZN(n91) );
  inv0d0 U130 ( .I(n72), .ZN(n39) );
  nd02d0 U131 ( .A1(n82), .A2(n83), .ZN(n111) );
  nd02d0 U132 ( .A1(n160), .A2(n86), .ZN(n112) );
  inv0d0 U133 ( .I(n53), .ZN(n35) );
  inv0d0 U134 ( .I(n64), .ZN(n37) );
  nd12d0 U135 ( .A1(n46), .A2(n45), .ZN(n104) );
  inv0d0 U136 ( .I(n58), .ZN(n60) );
  nd12d0 U137 ( .A1(n50), .A2(n49), .ZN(n105) );
  nd12d0 U138 ( .A1(n69), .A2(n68), .ZN(n109) );
  nd02d0 U139 ( .A1(A[9]), .A2(n26), .ZN(n86) );
  nd12d0 U140 ( .A1(n99), .A2(n98), .ZN(n114) );
  aoi21d1 U141 ( .B1(n57), .B2(n66), .A(n65), .ZN(n67) );
  aoi21d1 U142 ( .B1(n65), .B2(n74), .A(n73), .ZN(n75) );
  inv0d1 U143 ( .I(n84), .ZN(n82) );
  aoi21d1 U144 ( .B1(n47), .B2(n55), .A(n54), .ZN(n56) );
  aoi21d1 U145 ( .B1(n77), .B2(n96), .A(n95), .ZN(n97) );
  aoi21d1 U146 ( .B1(n160), .B2(n81), .A(n88), .ZN(n90) );
  inv0d1 U147 ( .I(n86), .ZN(n88) );
  inv0d1 U148 ( .I(n83), .ZN(n81) );
  nd12d0 U149 ( .A1(n94), .A2(n93), .ZN(n113) );
  inv0d1 U150 ( .I(n59), .ZN(n61) );
  xr02d1 U151 ( .A1(n158), .A2(n106), .Z(DIFF[3]) );
  ora21d1 U152 ( .B1(n48), .B2(n50), .A(n49), .Z(n158) );
  xn02d1 U153 ( .A1(n159), .A2(n108), .ZN(DIFF[5]) );
  aor21d1 U154 ( .B1(n57), .B2(n61), .A(n60), .Z(n159) );
  nd02d1 U155 ( .A1(A[4]), .A2(n21), .ZN(n58) );
  or02d1 U156 ( .A1(A[9]), .A2(n26), .Z(n160) );
  inv0d1 U157 ( .I(B[12]), .ZN(n29) );
  inv0d1 U158 ( .I(B[13]), .ZN(n30) );
  inv0d1 U159 ( .I(B[4]), .ZN(n21) );
  xn02d1 U160 ( .A1(B[15]), .A2(A[15]), .ZN(n115) );
  inv0d1 U161 ( .I(B[11]), .ZN(n28) );
  inv0d1 U162 ( .I(B[6]), .ZN(n23) );
  inv0d1 U163 ( .I(B[2]), .ZN(n19) );
  inv0d1 U164 ( .I(B[1]), .ZN(n18) );
  inv0d1 U165 ( .I(B[3]), .ZN(n20) );
  inv0d1 U166 ( .I(B[7]), .ZN(n24) );
  inv0d1 U167 ( .I(B[9]), .ZN(n26) );
  inv0d1 U168 ( .I(B[8]), .ZN(n25) );
  inv0d1 U169 ( .I(B[10]), .ZN(n27) );
  inv0d1 U170 ( .I(B[5]), .ZN(n22) );
  nd02d0 U171 ( .A1(A[5]), .A2(n22), .ZN(n63) );
endmodule


module PCI_FIFO_1_DW_fifoctl_s2_sf_0 ( clk_push, clk_pop, rst_n, push_req_n, 
        pop_req_n, we_n, push_empty, push_ae, push_hf, push_af, push_full, 
        push_error, pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, 
        wr_addr, rd_addr, push_word_count, pop_word_count, test, test_si1, 
        test_si2, test_se, test_so2, test_so1 );
  output [5:0] wr_addr;
  output [5:0] rd_addr;
  output [6:0] push_word_count;
  output [6:0] pop_word_count;
  input clk_push, clk_pop, rst_n, push_req_n, pop_req_n, test, test_si1,
         test_si2, test_se;
  output we_n, push_empty, push_ae, push_hf, push_af, push_full, push_error,
         pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, test_so2,
         test_so1;
  wire   rd_addr_gray_6_, rd_addr_gray_5_, rd_addr_gray_4_, rd_addr_gray_3_,
         rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_, wr_addr_gray_5_,
         wr_addr_gray_4_, wr_addr_gray_3_, wr_addr_gray_2_, wr_addr_gray_1_,
         wr_addr_gray_0_, SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68;

  PCI_FIFO_1_DW_FIFOCTL_IF_0 U2 ( .clk(clk_pop), .rst_n(rst_n), .init_n(1'b1), 
        .inc_req_n(pop_req_n), .other_addr_g({test_so2, wr_addr_gray_5_, 
        wr_addr_gray_4_, wr_addr_gray_3_, wr_addr_gray_2_, wr_addr_gray_1_, 
        wr_addr_gray_0_}), .word_count({SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41}), .empty(pop_empty), 
        .almost_empty(pop_ae), .half_full(pop_hf), .almost_full(pop_af), 
        .full(pop_full), .error(pop_error), .this_addr(rd_addr), .this_addr_g(
        {rd_addr_gray_6_, rd_addr_gray_5_, rd_addr_gray_4_, rd_addr_gray_3_, 
        rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_}), .next_word_count(
        {SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48}), .next_empty_n(SYNOPSYS_UNCONNECTED_49), 
        .next_full(SYNOPSYS_UNCONNECTED_50), .next_error(
        SYNOPSYS_UNCONNECTED_51), .test(test), .test_se(test_se), .test_si(
        test_si1), .test_so(test_so1) );
  PCI_FIFO_1_DW_FIFOCTL_IF_1 U1 ( .clk(clk_push), .rst_n(rst_n), .init_n(1'b1), 
        .inc_req_n(push_req_n), .other_addr_g({rd_addr_gray_6_, 
        rd_addr_gray_5_, rd_addr_gray_4_, rd_addr_gray_3_, rd_addr_gray_2_, 
        rd_addr_gray_1_, rd_addr_gray_0_}), .word_count({
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58}), .empty(push_empty), .almost_empty(push_ae), 
        .half_full(push_hf), .almost_full(push_af), .full(push_full), .error(
        push_error), .this_addr(wr_addr), .this_addr_g({test_so2, 
        wr_addr_gray_5_, wr_addr_gray_4_, wr_addr_gray_3_, wr_addr_gray_2_, 
        wr_addr_gray_1_, wr_addr_gray_0_}), .next_word_count({
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65}), .next_empty_n(SYNOPSYS_UNCONNECTED_66), 
        .next_full(SYNOPSYS_UNCONNECTED_67), .next_error(
        SYNOPSYS_UNCONNECTED_68), .test(test), .test_se(test_se), .test_si(
        test_si2) );
  or02d0 U6 ( .A1(push_full), .A2(push_req_n), .Z(we_n) );
endmodule


module PCI_FIFO_0_DW_fifoctl_s2_sf_0 ( clk_push, clk_pop, rst_n, push_req_n, 
        pop_req_n, we_n, push_empty, push_ae, push_hf, push_af, push_full, 
        push_error, pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, 
        wr_addr, rd_addr, push_word_count, pop_word_count, test, test_si1, 
        test_si2, test_se, test_so2, test_so1 );
  output [5:0] wr_addr;
  output [5:0] rd_addr;
  output [6:0] push_word_count;
  output [6:0] pop_word_count;
  input clk_push, clk_pop, rst_n, push_req_n, pop_req_n, test, test_si1,
         test_si2, test_se;
  output we_n, push_empty, push_ae, push_hf, push_af, push_full, push_error,
         pop_empty, pop_ae, pop_hf, pop_af, pop_full, pop_error, test_so2,
         test_so1;
  wire   rd_addr_gray_5_, rd_addr_gray_4_, rd_addr_gray_3_, rd_addr_gray_2_,
         rd_addr_gray_1_, rd_addr_gray_0_, wr_addr_gray_5_, wr_addr_gray_4_,
         wr_addr_gray_3_, wr_addr_gray_2_, wr_addr_gray_1_, wr_addr_gray_0_,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68;

  PCI_FIFO_0_DW_FIFOCTL_IF_0 U2 ( .clk(clk_pop), .rst_n(rst_n), .init_n(1'b1), 
        .inc_req_n(pop_req_n), .other_addr_g({test_so1, wr_addr_gray_5_, 
        wr_addr_gray_4_, wr_addr_gray_3_, wr_addr_gray_2_, wr_addr_gray_1_, 
        wr_addr_gray_0_}), .word_count({SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41}), .empty(pop_empty), 
        .almost_empty(pop_ae), .half_full(pop_hf), .almost_full(pop_af), 
        .full(pop_full), .error(pop_error), .this_addr(rd_addr), .this_addr_g(
        {test_so2, rd_addr_gray_5_, rd_addr_gray_4_, rd_addr_gray_3_, 
        rd_addr_gray_2_, rd_addr_gray_1_, rd_addr_gray_0_}), .next_word_count(
        {SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48}), .next_empty_n(SYNOPSYS_UNCONNECTED_49), 
        .next_full(SYNOPSYS_UNCONNECTED_50), .next_error(
        SYNOPSYS_UNCONNECTED_51), .test(test), .test_se(test_se), .test_si(
        test_si2) );
  PCI_FIFO_0_DW_FIFOCTL_IF_1 U1 ( .clk(clk_push), .rst_n(rst_n), .init_n(1'b1), 
        .inc_req_n(push_req_n), .other_addr_g({test_so2, rd_addr_gray_5_, 
        rd_addr_gray_4_, rd_addr_gray_3_, rd_addr_gray_2_, rd_addr_gray_1_, 
        rd_addr_gray_0_}), .word_count({SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58}), .empty(push_empty), 
        .almost_empty(push_ae), .half_full(push_hf), .almost_full(push_af), 
        .full(push_full), .error(push_error), .this_addr(wr_addr), 
        .this_addr_g({test_so1, wr_addr_gray_5_, wr_addr_gray_4_, 
        wr_addr_gray_3_, wr_addr_gray_2_, wr_addr_gray_1_, wr_addr_gray_0_}), 
        .next_word_count({SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65}), .next_empty_n(SYNOPSYS_UNCONNECTED_66), 
        .next_full(SYNOPSYS_UNCONNECTED_67), .next_error(
        SYNOPSYS_UNCONNECTED_68), .test(test), .test_se(test_se), .test_si(
        test_si1) );
  or02d0 U6 ( .A1(push_full), .A2(push_req_n), .Z(we_n) );
endmodule


module PCI_CORE_DW_mult_uns_3 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192;

  nr02d0 U17 ( .A1(n24), .A2(n16), .ZN(product[0]) );
  nr02d0 U18 ( .A1(n25), .A2(n16), .ZN(n33) );
  nr02d0 U19 ( .A1(n26), .A2(n16), .ZN(n34) );
  nr02d0 U20 ( .A1(n27), .A2(n16), .ZN(n35) );
  nr02d0 U21 ( .A1(n28), .A2(n16), .ZN(n36) );
  nr02d0 U22 ( .A1(n29), .A2(n16), .ZN(n37) );
  nr02d0 U23 ( .A1(n30), .A2(n16), .ZN(n38) );
  nr02d0 U24 ( .A1(n31), .A2(n16), .ZN(n39) );
  nr02d0 U25 ( .A1(n24), .A2(n17), .ZN(n40) );
  nr02d0 U26 ( .A1(n25), .A2(n17), .ZN(n41) );
  nr02d0 U27 ( .A1(n26), .A2(n17), .ZN(n42) );
  nr02d0 U28 ( .A1(n27), .A2(n17), .ZN(n43) );
  nr02d0 U29 ( .A1(n28), .A2(n17), .ZN(n44) );
  nr02d0 U30 ( .A1(n29), .A2(n17), .ZN(n45) );
  nr02d0 U31 ( .A1(n30), .A2(n17), .ZN(n46) );
  nr02d0 U32 ( .A1(n31), .A2(n17), .ZN(n47) );
  nr02d0 U33 ( .A1(n24), .A2(n18), .ZN(n48) );
  nr02d0 U34 ( .A1(n25), .A2(n18), .ZN(n49) );
  nr02d0 U35 ( .A1(n26), .A2(n18), .ZN(n50) );
  nr02d0 U36 ( .A1(n27), .A2(n18), .ZN(n51) );
  nr02d0 U37 ( .A1(n28), .A2(n18), .ZN(n52) );
  nr02d0 U38 ( .A1(n29), .A2(n18), .ZN(n53) );
  nr02d0 U39 ( .A1(n30), .A2(n18), .ZN(n54) );
  nr02d0 U40 ( .A1(n31), .A2(n18), .ZN(n55) );
  nr02d0 U41 ( .A1(n24), .A2(n19), .ZN(n56) );
  nr02d0 U42 ( .A1(n25), .A2(n19), .ZN(n57) );
  nr02d0 U43 ( .A1(n26), .A2(n19), .ZN(n58) );
  nr02d0 U44 ( .A1(n27), .A2(n19), .ZN(n59) );
  nr02d0 U45 ( .A1(n28), .A2(n19), .ZN(n60) );
  nr02d0 U46 ( .A1(n29), .A2(n19), .ZN(n61) );
  nr02d0 U47 ( .A1(n30), .A2(n19), .ZN(n62) );
  nr02d0 U48 ( .A1(n31), .A2(n19), .ZN(n63) );
  nr02d0 U49 ( .A1(n24), .A2(n20), .ZN(n64) );
  nr02d0 U50 ( .A1(n25), .A2(n20), .ZN(n65) );
  nr02d0 U51 ( .A1(n26), .A2(n20), .ZN(n66) );
  nr02d0 U52 ( .A1(n27), .A2(n20), .ZN(n67) );
  nr02d0 U53 ( .A1(n28), .A2(n20), .ZN(n68) );
  nr02d0 U54 ( .A1(n29), .A2(n20), .ZN(n69) );
  nr02d0 U55 ( .A1(n30), .A2(n20), .ZN(n70) );
  nr02d0 U56 ( .A1(n31), .A2(n20), .ZN(n71) );
  nr02d0 U57 ( .A1(n24), .A2(n21), .ZN(n72) );
  nr02d0 U58 ( .A1(n25), .A2(n21), .ZN(n73) );
  nr02d0 U59 ( .A1(n26), .A2(n21), .ZN(n74) );
  nr02d0 U60 ( .A1(n27), .A2(n21), .ZN(n75) );
  nr02d0 U61 ( .A1(n28), .A2(n21), .ZN(n76) );
  nr02d0 U62 ( .A1(n29), .A2(n21), .ZN(n77) );
  nr02d0 U63 ( .A1(n30), .A2(n21), .ZN(n78) );
  nr02d0 U64 ( .A1(n31), .A2(n21), .ZN(n79) );
  nr02d0 U65 ( .A1(n24), .A2(n22), .ZN(n80) );
  nr02d0 U66 ( .A1(n25), .A2(n22), .ZN(n81) );
  nr02d0 U67 ( .A1(n26), .A2(n22), .ZN(n82) );
  nr02d0 U68 ( .A1(n27), .A2(n22), .ZN(n83) );
  nr02d0 U69 ( .A1(n28), .A2(n22), .ZN(n84) );
  nr02d0 U70 ( .A1(n29), .A2(n22), .ZN(n85) );
  nr02d0 U71 ( .A1(n30), .A2(n22), .ZN(n86) );
  nr02d0 U72 ( .A1(n31), .A2(n22), .ZN(n87) );
  nr02d0 U73 ( .A1(n24), .A2(n23), .ZN(n88) );
  nr02d0 U74 ( .A1(n25), .A2(n23), .ZN(n89) );
  nr02d0 U75 ( .A1(n26), .A2(n23), .ZN(n90) );
  nr02d0 U76 ( .A1(n27), .A2(n23), .ZN(n91) );
  nr02d0 U77 ( .A1(n28), .A2(n23), .ZN(n92) );
  nr02d0 U78 ( .A1(n29), .A2(n23), .ZN(n93) );
  nr02d0 U79 ( .A1(n30), .A2(n23), .ZN(n94) );
  nr02d0 U80 ( .A1(n31), .A2(n23), .ZN(n95) );
  ah01d0 U81 ( .A(n34), .B(n41), .CO(n97), .S(n96) );
  ah01d0 U82 ( .A(n49), .B(n56), .CO(n99), .S(n98) );
  ad01d0 U83 ( .A(n35), .B(n42), .CI(n97), .CO(n101), .S(n100) );
  ah01d0 U84 ( .A(n57), .B(n64), .CO(n103), .S(n102) );
  ad01d0 U85 ( .A(n36), .B(n50), .CI(n43), .CO(n105), .S(n104) );
  ad01d0 U86 ( .A(n99), .B(n102), .CI(n104), .CO(n107), .S(n106) );
  ah01d0 U87 ( .A(n65), .B(n72), .CO(n109), .S(n108) );
  ad01d0 U88 ( .A(n37), .B(n58), .CI(n51), .CO(n111), .S(n110) );
  ad01d0 U89 ( .A(n44), .B(n103), .CI(n108), .CO(n113), .S(n112) );
  ad01d0 U90 ( .A(n105), .B(n110), .CI(n112), .CO(n115), .S(n114) );
  ah01d0 U91 ( .A(n73), .B(n80), .CO(n117), .S(n116) );
  ad01d0 U92 ( .A(n38), .B(n66), .CI(n45), .CO(n119), .S(n118) );
  ad01d0 U93 ( .A(n52), .B(n59), .CI(n109), .CO(n121), .S(n120) );
  ad01d0 U94 ( .A(n116), .B(n111), .CI(n118), .CO(n123), .S(n122) );
  ad01d0 U95 ( .A(n113), .B(n120), .CI(n122), .CO(n125), .S(n124) );
  ah01d0 U96 ( .A(n81), .B(n88), .CO(n127), .S(n126) );
  ad01d0 U97 ( .A(n39), .B(n74), .CI(n46), .CO(n129), .S(n128) );
  ad01d0 U98 ( .A(n53), .B(n67), .CI(n60), .CO(n131), .S(n130) );
  ad01d0 U99 ( .A(n117), .B(n126), .CI(n119), .CO(n133), .S(n132) );
  ad01d0 U100 ( .A(n130), .B(n128), .CI(n121), .CO(n135), .S(n134) );
  ad01d0 U101 ( .A(n132), .B(n123), .CI(n134), .CO(n137), .S(n136) );
  ah01d0 U102 ( .A(n82), .B(n89), .CO(n139), .S(n138) );
  ad01d0 U103 ( .A(n68), .B(n75), .CI(n47), .CO(n141), .S(n140) );
  ad01d0 U104 ( .A(n54), .B(n61), .CI(n127), .CO(n143), .S(n142) );
  ad01d0 U105 ( .A(n138), .B(n129), .CI(n131), .CO(n145), .S(n144) );
  ad01d0 U106 ( .A(n140), .B(n142), .CI(n133), .CO(n147), .S(n146) );
  ad01d0 U107 ( .A(n144), .B(n135), .CI(n146), .CO(n149), .S(n148) );
  ad01d0 U108 ( .A(n55), .B(n90), .CI(n83), .CO(n151), .S(n150) );
  ad01d0 U109 ( .A(n76), .B(n69), .CI(n62), .CO(n153), .S(n152) );
  ad01d0 U110 ( .A(n139), .B(n141), .CI(n152), .CO(n155), .S(n154) );
  ad01d0 U111 ( .A(n150), .B(n143), .CI(n145), .CO(n157), .S(n156) );
  ad01d0 U112 ( .A(n154), .B(n147), .CI(n156), .CO(n159), .S(n158) );
  ad01d0 U113 ( .A(n63), .B(n91), .CI(n84), .CO(n161), .S(n160) );
  ad01d0 U114 ( .A(n70), .B(n77), .CI(n151), .CO(n163), .S(n162) );
  ad01d0 U115 ( .A(n153), .B(n160), .CI(n162), .CO(n165), .S(n164) );
  ad01d0 U116 ( .A(n155), .B(n157), .CI(n164), .CO(n167), .S(n166) );
  ad01d0 U117 ( .A(n71), .B(n92), .CI(n85), .CO(n169), .S(n168) );
  ad01d0 U118 ( .A(n78), .B(n161), .CI(n168), .CO(n171), .S(n170) );
  ad01d0 U119 ( .A(n163), .B(n170), .CI(n165), .CO(n173), .S(n172) );
  ad01d0 U120 ( .A(n79), .B(n93), .CI(n86), .CO(n175), .S(n174) );
  ad01d0 U121 ( .A(n169), .B(n174), .CI(n171), .CO(n177), .S(n176) );
  ad01d0 U122 ( .A(n87), .B(n94), .CI(n175), .CO(n179), .S(n178) );
  ah01d0 U123 ( .A(n40), .B(n33), .CO(n180), .S(product[1]) );
  ad01d0 U124 ( .A(n48), .B(n180), .CI(n96), .CO(n181), .S(product[2]) );
  ad01d0 U125 ( .A(n98), .B(n181), .CI(n100), .CO(n182), .S(product[3]) );
  ad01d0 U126 ( .A(n101), .B(n106), .CI(n182), .CO(n183), .S(product[4]) );
  ad01d0 U127 ( .A(n107), .B(n114), .CI(n183), .CO(n184), .S(product[5]) );
  ad01d0 U128 ( .A(n115), .B(n124), .CI(n184), .CO(n185), .S(product[6]) );
  ad01d0 U129 ( .A(n125), .B(n136), .CI(n185), .CO(n186), .S(product[7]) );
  ad01d0 U130 ( .A(n137), .B(n148), .CI(n186), .CO(n187), .S(product[8]) );
  ad01d0 U131 ( .A(n149), .B(n158), .CI(n187), .CO(n188), .S(product[9]) );
  ad01d0 U132 ( .A(n159), .B(n166), .CI(n188), .CO(n189), .S(product[10]) );
  ad01d0 U133 ( .A(n167), .B(n172), .CI(n189), .CO(n190), .S(product[11]) );
  ad01d0 U134 ( .A(n176), .B(n173), .CI(n190), .CO(n191), .S(product[12]) );
  ad01d0 U135 ( .A(n178), .B(n177), .CI(n191), .CO(n192), .S(product[13]) );
  ad01d0 U136 ( .A(n95), .B(n179), .CI(n192), .CO(product[15]), .S(product[14]) );
  inv0d1 U140 ( .I(a[4]), .ZN(n20) );
  inv0d1 U141 ( .I(a[3]), .ZN(n19) );
  inv0d1 U142 ( .I(a[0]), .ZN(n16) );
  inv0d1 U143 ( .I(a[2]), .ZN(n18) );
  inv0d1 U144 ( .I(a[1]), .ZN(n17) );
  inv0d1 U145 ( .I(a[5]), .ZN(n21) );
  inv0d1 U146 ( .I(a[6]), .ZN(n22) );
  inv0d1 U147 ( .I(a[7]), .ZN(n23) );
  inv0d1 U148 ( .I(b[1]), .ZN(n25) );
  inv0d1 U149 ( .I(b[0]), .ZN(n24) );
  inv0d1 U150 ( .I(b[2]), .ZN(n26) );
  inv0d1 U151 ( .I(b[3]), .ZN(n27) );
  inv0d1 U152 ( .I(b[4]), .ZN(n28) );
  inv0d1 U153 ( .I(b[5]), .ZN(n29) );
  inv0d1 U154 ( .I(b[6]), .ZN(n30) );
  inv0d1 U155 ( .I(b[7]), .ZN(n31) );
endmodule


module PCI_CORE_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192;

  nr02d0 U17 ( .A1(n24), .A2(n16), .ZN(product[0]) );
  nr02d0 U18 ( .A1(n25), .A2(n16), .ZN(n33) );
  nr02d0 U19 ( .A1(n26), .A2(n16), .ZN(n34) );
  nr02d0 U20 ( .A1(n27), .A2(n16), .ZN(n35) );
  nr02d0 U21 ( .A1(n28), .A2(n16), .ZN(n36) );
  nr02d0 U22 ( .A1(n29), .A2(n16), .ZN(n37) );
  nr02d0 U23 ( .A1(n30), .A2(n16), .ZN(n38) );
  nr02d0 U24 ( .A1(n31), .A2(n16), .ZN(n39) );
  nr02d0 U25 ( .A1(n24), .A2(n17), .ZN(n40) );
  nr02d0 U26 ( .A1(n25), .A2(n17), .ZN(n41) );
  nr02d0 U27 ( .A1(n26), .A2(n17), .ZN(n42) );
  nr02d0 U28 ( .A1(n27), .A2(n17), .ZN(n43) );
  nr02d0 U29 ( .A1(n28), .A2(n17), .ZN(n44) );
  nr02d0 U30 ( .A1(n29), .A2(n17), .ZN(n45) );
  nr02d0 U31 ( .A1(n30), .A2(n17), .ZN(n46) );
  nr02d0 U32 ( .A1(n31), .A2(n17), .ZN(n47) );
  nr02d0 U33 ( .A1(n24), .A2(n18), .ZN(n48) );
  nr02d0 U34 ( .A1(n25), .A2(n18), .ZN(n49) );
  nr02d0 U35 ( .A1(n26), .A2(n18), .ZN(n50) );
  nr02d0 U36 ( .A1(n27), .A2(n18), .ZN(n51) );
  nr02d0 U37 ( .A1(n28), .A2(n18), .ZN(n52) );
  nr02d0 U38 ( .A1(n29), .A2(n18), .ZN(n53) );
  nr02d0 U39 ( .A1(n30), .A2(n18), .ZN(n54) );
  nr02d0 U40 ( .A1(n31), .A2(n18), .ZN(n55) );
  nr02d0 U41 ( .A1(n24), .A2(n19), .ZN(n56) );
  nr02d0 U42 ( .A1(n25), .A2(n19), .ZN(n57) );
  nr02d0 U43 ( .A1(n26), .A2(n19), .ZN(n58) );
  nr02d0 U44 ( .A1(n27), .A2(n19), .ZN(n59) );
  nr02d0 U45 ( .A1(n28), .A2(n19), .ZN(n60) );
  nr02d0 U46 ( .A1(n29), .A2(n19), .ZN(n61) );
  nr02d0 U47 ( .A1(n30), .A2(n19), .ZN(n62) );
  nr02d0 U48 ( .A1(n31), .A2(n19), .ZN(n63) );
  nr02d0 U49 ( .A1(n24), .A2(n20), .ZN(n64) );
  nr02d0 U50 ( .A1(n25), .A2(n20), .ZN(n65) );
  nr02d0 U51 ( .A1(n26), .A2(n20), .ZN(n66) );
  nr02d0 U52 ( .A1(n27), .A2(n20), .ZN(n67) );
  nr02d0 U53 ( .A1(n28), .A2(n20), .ZN(n68) );
  nr02d0 U54 ( .A1(n29), .A2(n20), .ZN(n69) );
  nr02d0 U55 ( .A1(n30), .A2(n20), .ZN(n70) );
  nr02d0 U56 ( .A1(n31), .A2(n20), .ZN(n71) );
  nr02d0 U57 ( .A1(n24), .A2(n21), .ZN(n72) );
  nr02d0 U58 ( .A1(n25), .A2(n21), .ZN(n73) );
  nr02d0 U59 ( .A1(n26), .A2(n21), .ZN(n74) );
  nr02d0 U60 ( .A1(n27), .A2(n21), .ZN(n75) );
  nr02d0 U61 ( .A1(n28), .A2(n21), .ZN(n76) );
  nr02d0 U62 ( .A1(n29), .A2(n21), .ZN(n77) );
  nr02d0 U63 ( .A1(n30), .A2(n21), .ZN(n78) );
  nr02d0 U64 ( .A1(n31), .A2(n21), .ZN(n79) );
  nr02d0 U65 ( .A1(n24), .A2(n22), .ZN(n80) );
  nr02d0 U66 ( .A1(n25), .A2(n22), .ZN(n81) );
  nr02d0 U67 ( .A1(n26), .A2(n22), .ZN(n82) );
  nr02d0 U68 ( .A1(n27), .A2(n22), .ZN(n83) );
  nr02d0 U69 ( .A1(n28), .A2(n22), .ZN(n84) );
  nr02d0 U70 ( .A1(n29), .A2(n22), .ZN(n85) );
  nr02d0 U71 ( .A1(n30), .A2(n22), .ZN(n86) );
  nr02d0 U72 ( .A1(n31), .A2(n22), .ZN(n87) );
  nr02d0 U73 ( .A1(n24), .A2(n23), .ZN(n88) );
  nr02d0 U74 ( .A1(n25), .A2(n23), .ZN(n89) );
  nr02d0 U75 ( .A1(n26), .A2(n23), .ZN(n90) );
  nr02d0 U76 ( .A1(n27), .A2(n23), .ZN(n91) );
  nr02d0 U77 ( .A1(n28), .A2(n23), .ZN(n92) );
  nr02d0 U78 ( .A1(n29), .A2(n23), .ZN(n93) );
  nr02d0 U79 ( .A1(n30), .A2(n23), .ZN(n94) );
  nr02d0 U80 ( .A1(n31), .A2(n23), .ZN(n95) );
  ah01d0 U81 ( .A(n34), .B(n41), .CO(n97), .S(n96) );
  ah01d0 U82 ( .A(n49), .B(n56), .CO(n99), .S(n98) );
  ad01d0 U83 ( .A(n35), .B(n42), .CI(n97), .CO(n101), .S(n100) );
  ah01d0 U84 ( .A(n57), .B(n64), .CO(n103), .S(n102) );
  ad01d0 U85 ( .A(n36), .B(n50), .CI(n43), .CO(n105), .S(n104) );
  ad01d0 U86 ( .A(n99), .B(n102), .CI(n104), .CO(n107), .S(n106) );
  ah01d0 U87 ( .A(n65), .B(n72), .CO(n109), .S(n108) );
  ad01d0 U88 ( .A(n37), .B(n58), .CI(n51), .CO(n111), .S(n110) );
  ad01d0 U89 ( .A(n44), .B(n103), .CI(n108), .CO(n113), .S(n112) );
  ad01d0 U90 ( .A(n105), .B(n110), .CI(n112), .CO(n115), .S(n114) );
  ah01d0 U91 ( .A(n73), .B(n80), .CO(n117), .S(n116) );
  ad01d0 U92 ( .A(n38), .B(n66), .CI(n45), .CO(n119), .S(n118) );
  ad01d0 U93 ( .A(n52), .B(n59), .CI(n109), .CO(n121), .S(n120) );
  ad01d0 U94 ( .A(n116), .B(n111), .CI(n118), .CO(n123), .S(n122) );
  ad01d0 U95 ( .A(n113), .B(n120), .CI(n122), .CO(n125), .S(n124) );
  ah01d0 U96 ( .A(n81), .B(n88), .CO(n127), .S(n126) );
  ad01d0 U97 ( .A(n39), .B(n74), .CI(n46), .CO(n129), .S(n128) );
  ad01d0 U98 ( .A(n53), .B(n67), .CI(n60), .CO(n131), .S(n130) );
  ad01d0 U99 ( .A(n117), .B(n126), .CI(n119), .CO(n133), .S(n132) );
  ad01d0 U100 ( .A(n130), .B(n128), .CI(n121), .CO(n135), .S(n134) );
  ad01d0 U101 ( .A(n132), .B(n123), .CI(n134), .CO(n137), .S(n136) );
  ah01d0 U102 ( .A(n82), .B(n89), .CO(n139), .S(n138) );
  ad01d0 U103 ( .A(n68), .B(n75), .CI(n47), .CO(n141), .S(n140) );
  ad01d0 U104 ( .A(n54), .B(n61), .CI(n127), .CO(n143), .S(n142) );
  ad01d0 U105 ( .A(n138), .B(n129), .CI(n131), .CO(n145), .S(n144) );
  ad01d0 U106 ( .A(n140), .B(n142), .CI(n133), .CO(n147), .S(n146) );
  ad01d0 U107 ( .A(n144), .B(n135), .CI(n146), .CO(n149), .S(n148) );
  ad01d0 U108 ( .A(n55), .B(n90), .CI(n83), .CO(n151), .S(n150) );
  ad01d0 U109 ( .A(n76), .B(n69), .CI(n62), .CO(n153), .S(n152) );
  ad01d0 U110 ( .A(n139), .B(n141), .CI(n152), .CO(n155), .S(n154) );
  ad01d0 U111 ( .A(n150), .B(n143), .CI(n145), .CO(n157), .S(n156) );
  ad01d0 U112 ( .A(n154), .B(n147), .CI(n156), .CO(n159), .S(n158) );
  ad01d0 U113 ( .A(n63), .B(n91), .CI(n84), .CO(n161), .S(n160) );
  ad01d0 U114 ( .A(n70), .B(n77), .CI(n151), .CO(n163), .S(n162) );
  ad01d0 U115 ( .A(n153), .B(n160), .CI(n162), .CO(n165), .S(n164) );
  ad01d0 U116 ( .A(n155), .B(n157), .CI(n164), .CO(n167), .S(n166) );
  ad01d0 U117 ( .A(n71), .B(n92), .CI(n85), .CO(n169), .S(n168) );
  ad01d0 U118 ( .A(n78), .B(n161), .CI(n168), .CO(n171), .S(n170) );
  ad01d0 U119 ( .A(n163), .B(n170), .CI(n165), .CO(n173), .S(n172) );
  ad01d0 U120 ( .A(n79), .B(n93), .CI(n86), .CO(n175), .S(n174) );
  ad01d0 U121 ( .A(n169), .B(n174), .CI(n171), .CO(n177), .S(n176) );
  ad01d0 U122 ( .A(n87), .B(n94), .CI(n175), .CO(n179), .S(n178) );
  ah01d0 U123 ( .A(n40), .B(n33), .CO(n180), .S(product[1]) );
  ad01d0 U124 ( .A(n48), .B(n180), .CI(n96), .CO(n181), .S(product[2]) );
  ad01d0 U125 ( .A(n98), .B(n181), .CI(n100), .CO(n182), .S(product[3]) );
  ad01d0 U126 ( .A(n101), .B(n106), .CI(n182), .CO(n183), .S(product[4]) );
  ad01d0 U127 ( .A(n107), .B(n114), .CI(n183), .CO(n184), .S(product[5]) );
  ad01d0 U128 ( .A(n115), .B(n124), .CI(n184), .CO(n185), .S(product[6]) );
  ad01d0 U129 ( .A(n125), .B(n136), .CI(n185), .CO(n186), .S(product[7]) );
  ad01d0 U130 ( .A(n137), .B(n148), .CI(n186), .CO(n187), .S(product[8]) );
  ad01d0 U131 ( .A(n149), .B(n158), .CI(n187), .CO(n188), .S(product[9]) );
  ad01d0 U132 ( .A(n159), .B(n166), .CI(n188), .CO(n189), .S(product[10]) );
  ad01d0 U133 ( .A(n167), .B(n172), .CI(n189), .CO(n190), .S(product[11]) );
  ad01d0 U134 ( .A(n176), .B(n173), .CI(n190), .CO(n191), .S(product[12]) );
  ad01d0 U135 ( .A(n178), .B(n177), .CI(n191), .CO(n192), .S(product[13]) );
  ad01d0 U136 ( .A(n95), .B(n179), .CI(n192), .CO(product[15]), .S(product[14]) );
  inv0d1 U140 ( .I(a[4]), .ZN(n20) );
  inv0d1 U141 ( .I(a[3]), .ZN(n19) );
  inv0d1 U142 ( .I(a[0]), .ZN(n16) );
  inv0d1 U143 ( .I(a[2]), .ZN(n18) );
  inv0d1 U144 ( .I(a[1]), .ZN(n17) );
  inv0d1 U145 ( .I(a[5]), .ZN(n21) );
  inv0d1 U146 ( .I(a[6]), .ZN(n22) );
  inv0d1 U147 ( .I(a[7]), .ZN(n23) );
  inv0d1 U148 ( .I(b[1]), .ZN(n25) );
  inv0d1 U149 ( .I(b[0]), .ZN(n24) );
  inv0d1 U150 ( .I(b[2]), .ZN(n26) );
  inv0d1 U151 ( .I(b[3]), .ZN(n27) );
  inv0d1 U152 ( .I(b[4]), .ZN(n28) );
  inv0d1 U153 ( .I(b[5]), .ZN(n29) );
  inv0d1 U154 ( .I(b[6]), .ZN(n30) );
  inv0d1 U155 ( .I(b[7]), .ZN(n31) );
endmodule


module PCI_CORE_DW_mult_uns_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192;

  nr02d0 U17 ( .A1(n24), .A2(n16), .ZN(product[0]) );
  nr02d0 U18 ( .A1(n25), .A2(n16), .ZN(n33) );
  nr02d0 U19 ( .A1(n26), .A2(n16), .ZN(n34) );
  nr02d0 U20 ( .A1(n27), .A2(n16), .ZN(n35) );
  nr02d0 U21 ( .A1(n28), .A2(n16), .ZN(n36) );
  nr02d0 U22 ( .A1(n29), .A2(n16), .ZN(n37) );
  nr02d0 U23 ( .A1(n30), .A2(n16), .ZN(n38) );
  nr02d0 U24 ( .A1(n31), .A2(n16), .ZN(n39) );
  nr02d0 U25 ( .A1(n24), .A2(n17), .ZN(n40) );
  nr02d0 U26 ( .A1(n25), .A2(n17), .ZN(n41) );
  nr02d0 U27 ( .A1(n26), .A2(n17), .ZN(n42) );
  nr02d0 U28 ( .A1(n27), .A2(n17), .ZN(n43) );
  nr02d0 U29 ( .A1(n28), .A2(n17), .ZN(n44) );
  nr02d0 U30 ( .A1(n29), .A2(n17), .ZN(n45) );
  nr02d0 U31 ( .A1(n30), .A2(n17), .ZN(n46) );
  nr02d0 U32 ( .A1(n31), .A2(n17), .ZN(n47) );
  nr02d0 U33 ( .A1(n24), .A2(n18), .ZN(n48) );
  nr02d0 U34 ( .A1(n25), .A2(n18), .ZN(n49) );
  nr02d0 U35 ( .A1(n26), .A2(n18), .ZN(n50) );
  nr02d0 U36 ( .A1(n27), .A2(n18), .ZN(n51) );
  nr02d0 U37 ( .A1(n28), .A2(n18), .ZN(n52) );
  nr02d0 U38 ( .A1(n29), .A2(n18), .ZN(n53) );
  nr02d0 U39 ( .A1(n30), .A2(n18), .ZN(n54) );
  nr02d0 U40 ( .A1(n31), .A2(n18), .ZN(n55) );
  nr02d0 U41 ( .A1(n24), .A2(n19), .ZN(n56) );
  nr02d0 U42 ( .A1(n25), .A2(n19), .ZN(n57) );
  nr02d0 U43 ( .A1(n26), .A2(n19), .ZN(n58) );
  nr02d0 U44 ( .A1(n27), .A2(n19), .ZN(n59) );
  nr02d0 U45 ( .A1(n28), .A2(n19), .ZN(n60) );
  nr02d0 U46 ( .A1(n29), .A2(n19), .ZN(n61) );
  nr02d0 U47 ( .A1(n30), .A2(n19), .ZN(n62) );
  nr02d0 U48 ( .A1(n31), .A2(n19), .ZN(n63) );
  nr02d0 U49 ( .A1(n24), .A2(n20), .ZN(n64) );
  nr02d0 U50 ( .A1(n25), .A2(n20), .ZN(n65) );
  nr02d0 U51 ( .A1(n26), .A2(n20), .ZN(n66) );
  nr02d0 U52 ( .A1(n27), .A2(n20), .ZN(n67) );
  nr02d0 U53 ( .A1(n28), .A2(n20), .ZN(n68) );
  nr02d0 U54 ( .A1(n29), .A2(n20), .ZN(n69) );
  nr02d0 U55 ( .A1(n30), .A2(n20), .ZN(n70) );
  nr02d0 U56 ( .A1(n31), .A2(n20), .ZN(n71) );
  nr02d0 U57 ( .A1(n24), .A2(n21), .ZN(n72) );
  nr02d0 U58 ( .A1(n25), .A2(n21), .ZN(n73) );
  nr02d0 U59 ( .A1(n26), .A2(n21), .ZN(n74) );
  nr02d0 U60 ( .A1(n27), .A2(n21), .ZN(n75) );
  nr02d0 U61 ( .A1(n28), .A2(n21), .ZN(n76) );
  nr02d0 U62 ( .A1(n29), .A2(n21), .ZN(n77) );
  nr02d0 U63 ( .A1(n30), .A2(n21), .ZN(n78) );
  nr02d0 U64 ( .A1(n31), .A2(n21), .ZN(n79) );
  nr02d0 U65 ( .A1(n24), .A2(n22), .ZN(n80) );
  nr02d0 U66 ( .A1(n25), .A2(n22), .ZN(n81) );
  nr02d0 U67 ( .A1(n26), .A2(n22), .ZN(n82) );
  nr02d0 U68 ( .A1(n27), .A2(n22), .ZN(n83) );
  nr02d0 U69 ( .A1(n28), .A2(n22), .ZN(n84) );
  nr02d0 U70 ( .A1(n29), .A2(n22), .ZN(n85) );
  nr02d0 U71 ( .A1(n30), .A2(n22), .ZN(n86) );
  nr02d0 U72 ( .A1(n31), .A2(n22), .ZN(n87) );
  nr02d0 U73 ( .A1(n24), .A2(n23), .ZN(n88) );
  nr02d0 U74 ( .A1(n25), .A2(n23), .ZN(n89) );
  nr02d0 U75 ( .A1(n26), .A2(n23), .ZN(n90) );
  nr02d0 U76 ( .A1(n27), .A2(n23), .ZN(n91) );
  nr02d0 U77 ( .A1(n28), .A2(n23), .ZN(n92) );
  nr02d0 U78 ( .A1(n29), .A2(n23), .ZN(n93) );
  nr02d0 U79 ( .A1(n30), .A2(n23), .ZN(n94) );
  nr02d0 U80 ( .A1(n31), .A2(n23), .ZN(n95) );
  ah01d0 U81 ( .A(n34), .B(n41), .CO(n97), .S(n96) );
  ah01d0 U82 ( .A(n49), .B(n56), .CO(n99), .S(n98) );
  ad01d0 U83 ( .A(n35), .B(n42), .CI(n97), .CO(n101), .S(n100) );
  ah01d0 U84 ( .A(n57), .B(n64), .CO(n103), .S(n102) );
  ad01d0 U85 ( .A(n36), .B(n50), .CI(n43), .CO(n105), .S(n104) );
  ad01d0 U86 ( .A(n99), .B(n102), .CI(n104), .CO(n107), .S(n106) );
  ah01d0 U87 ( .A(n65), .B(n72), .CO(n109), .S(n108) );
  ad01d0 U88 ( .A(n37), .B(n58), .CI(n51), .CO(n111), .S(n110) );
  ad01d0 U89 ( .A(n44), .B(n103), .CI(n108), .CO(n113), .S(n112) );
  ad01d0 U90 ( .A(n105), .B(n110), .CI(n112), .CO(n115), .S(n114) );
  ah01d0 U91 ( .A(n73), .B(n80), .CO(n117), .S(n116) );
  ad01d0 U92 ( .A(n38), .B(n66), .CI(n45), .CO(n119), .S(n118) );
  ad01d0 U93 ( .A(n52), .B(n59), .CI(n109), .CO(n121), .S(n120) );
  ad01d0 U94 ( .A(n116), .B(n111), .CI(n118), .CO(n123), .S(n122) );
  ad01d0 U95 ( .A(n113), .B(n120), .CI(n122), .CO(n125), .S(n124) );
  ah01d0 U96 ( .A(n81), .B(n88), .CO(n127), .S(n126) );
  ad01d0 U97 ( .A(n39), .B(n74), .CI(n46), .CO(n129), .S(n128) );
  ad01d0 U98 ( .A(n53), .B(n67), .CI(n60), .CO(n131), .S(n130) );
  ad01d0 U99 ( .A(n117), .B(n126), .CI(n119), .CO(n133), .S(n132) );
  ad01d0 U100 ( .A(n130), .B(n128), .CI(n121), .CO(n135), .S(n134) );
  ad01d0 U101 ( .A(n132), .B(n123), .CI(n134), .CO(n137), .S(n136) );
  ah01d0 U102 ( .A(n82), .B(n89), .CO(n139), .S(n138) );
  ad01d0 U103 ( .A(n68), .B(n75), .CI(n47), .CO(n141), .S(n140) );
  ad01d0 U104 ( .A(n54), .B(n61), .CI(n127), .CO(n143), .S(n142) );
  ad01d0 U105 ( .A(n138), .B(n129), .CI(n131), .CO(n145), .S(n144) );
  ad01d0 U106 ( .A(n140), .B(n142), .CI(n133), .CO(n147), .S(n146) );
  ad01d0 U107 ( .A(n144), .B(n135), .CI(n146), .CO(n149), .S(n148) );
  ad01d0 U108 ( .A(n55), .B(n90), .CI(n83), .CO(n151), .S(n150) );
  ad01d0 U109 ( .A(n76), .B(n69), .CI(n62), .CO(n153), .S(n152) );
  ad01d0 U110 ( .A(n139), .B(n141), .CI(n152), .CO(n155), .S(n154) );
  ad01d0 U111 ( .A(n150), .B(n143), .CI(n145), .CO(n157), .S(n156) );
  ad01d0 U112 ( .A(n154), .B(n147), .CI(n156), .CO(n159), .S(n158) );
  ad01d0 U113 ( .A(n63), .B(n91), .CI(n84), .CO(n161), .S(n160) );
  ad01d0 U114 ( .A(n70), .B(n77), .CI(n151), .CO(n163), .S(n162) );
  ad01d0 U115 ( .A(n153), .B(n160), .CI(n162), .CO(n165), .S(n164) );
  ad01d0 U116 ( .A(n155), .B(n157), .CI(n164), .CO(n167), .S(n166) );
  ad01d0 U117 ( .A(n71), .B(n92), .CI(n85), .CO(n169), .S(n168) );
  ad01d0 U118 ( .A(n78), .B(n161), .CI(n168), .CO(n171), .S(n170) );
  ad01d0 U119 ( .A(n163), .B(n170), .CI(n165), .CO(n173), .S(n172) );
  ad01d0 U120 ( .A(n79), .B(n93), .CI(n86), .CO(n175), .S(n174) );
  ad01d0 U121 ( .A(n169), .B(n174), .CI(n171), .CO(n177), .S(n176) );
  ad01d0 U122 ( .A(n87), .B(n94), .CI(n175), .CO(n179), .S(n178) );
  ah01d0 U123 ( .A(n40), .B(n33), .CO(n180), .S(product[1]) );
  ad01d0 U124 ( .A(n48), .B(n180), .CI(n96), .CO(n181), .S(product[2]) );
  ad01d0 U125 ( .A(n98), .B(n181), .CI(n100), .CO(n182), .S(product[3]) );
  ad01d0 U126 ( .A(n101), .B(n106), .CI(n182), .CO(n183), .S(product[4]) );
  ad01d0 U127 ( .A(n107), .B(n114), .CI(n183), .CO(n184), .S(product[5]) );
  ad01d0 U128 ( .A(n115), .B(n124), .CI(n184), .CO(n185), .S(product[6]) );
  ad01d0 U129 ( .A(n125), .B(n136), .CI(n185), .CO(n186), .S(product[7]) );
  ad01d0 U130 ( .A(n137), .B(n148), .CI(n186), .CO(n187), .S(product[8]) );
  ad01d0 U131 ( .A(n149), .B(n158), .CI(n187), .CO(n188), .S(product[9]) );
  ad01d0 U132 ( .A(n159), .B(n166), .CI(n188), .CO(n189), .S(product[10]) );
  ad01d0 U133 ( .A(n167), .B(n172), .CI(n189), .CO(n190), .S(product[11]) );
  ad01d0 U134 ( .A(n176), .B(n173), .CI(n190), .CO(n191), .S(product[12]) );
  ad01d0 U135 ( .A(n178), .B(n177), .CI(n191), .CO(n192), .S(product[13]) );
  ad01d0 U136 ( .A(n95), .B(n179), .CI(n192), .CO(product[15]), .S(product[14]) );
  inv0d1 U140 ( .I(a[4]), .ZN(n20) );
  inv0d1 U141 ( .I(a[3]), .ZN(n19) );
  inv0d1 U142 ( .I(a[0]), .ZN(n16) );
  inv0d1 U143 ( .I(a[2]), .ZN(n18) );
  inv0d1 U144 ( .I(a[1]), .ZN(n17) );
  inv0d1 U145 ( .I(a[5]), .ZN(n21) );
  inv0d1 U146 ( .I(a[6]), .ZN(n22) );
  inv0d1 U147 ( .I(a[7]), .ZN(n23) );
  inv0d1 U148 ( .I(b[1]), .ZN(n25) );
  inv0d1 U149 ( .I(b[0]), .ZN(n24) );
  inv0d1 U150 ( .I(b[2]), .ZN(n26) );
  inv0d1 U151 ( .I(b[3]), .ZN(n27) );
  inv0d1 U152 ( .I(b[4]), .ZN(n28) );
  inv0d1 U153 ( .I(b[5]), .ZN(n29) );
  inv0d1 U154 ( .I(b[6]), .ZN(n30) );
  inv0d1 U155 ( .I(b[7]), .ZN(n31) );
endmodule


module PCI_CORE_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192;

  nr02d0 U17 ( .A1(n24), .A2(n16), .ZN(product[0]) );
  nr02d0 U18 ( .A1(n25), .A2(n16), .ZN(n33) );
  nr02d0 U19 ( .A1(n26), .A2(n16), .ZN(n34) );
  nr02d0 U20 ( .A1(n27), .A2(n16), .ZN(n35) );
  nr02d0 U21 ( .A1(n28), .A2(n16), .ZN(n36) );
  nr02d0 U22 ( .A1(n29), .A2(n16), .ZN(n37) );
  nr02d0 U23 ( .A1(n30), .A2(n16), .ZN(n38) );
  nr02d0 U24 ( .A1(n31), .A2(n16), .ZN(n39) );
  nr02d0 U25 ( .A1(n24), .A2(n17), .ZN(n40) );
  nr02d0 U26 ( .A1(n25), .A2(n17), .ZN(n41) );
  nr02d0 U27 ( .A1(n26), .A2(n17), .ZN(n42) );
  nr02d0 U28 ( .A1(n27), .A2(n17), .ZN(n43) );
  nr02d0 U29 ( .A1(n28), .A2(n17), .ZN(n44) );
  nr02d0 U30 ( .A1(n29), .A2(n17), .ZN(n45) );
  nr02d0 U31 ( .A1(n30), .A2(n17), .ZN(n46) );
  nr02d0 U32 ( .A1(n31), .A2(n17), .ZN(n47) );
  nr02d0 U33 ( .A1(n24), .A2(n18), .ZN(n48) );
  nr02d0 U34 ( .A1(n25), .A2(n18), .ZN(n49) );
  nr02d0 U35 ( .A1(n26), .A2(n18), .ZN(n50) );
  nr02d0 U36 ( .A1(n27), .A2(n18), .ZN(n51) );
  nr02d0 U37 ( .A1(n28), .A2(n18), .ZN(n52) );
  nr02d0 U38 ( .A1(n29), .A2(n18), .ZN(n53) );
  nr02d0 U39 ( .A1(n30), .A2(n18), .ZN(n54) );
  nr02d0 U40 ( .A1(n31), .A2(n18), .ZN(n55) );
  nr02d0 U41 ( .A1(n24), .A2(n19), .ZN(n56) );
  nr02d0 U42 ( .A1(n25), .A2(n19), .ZN(n57) );
  nr02d0 U43 ( .A1(n26), .A2(n19), .ZN(n58) );
  nr02d0 U44 ( .A1(n27), .A2(n19), .ZN(n59) );
  nr02d0 U45 ( .A1(n28), .A2(n19), .ZN(n60) );
  nr02d0 U46 ( .A1(n29), .A2(n19), .ZN(n61) );
  nr02d0 U47 ( .A1(n30), .A2(n19), .ZN(n62) );
  nr02d0 U48 ( .A1(n31), .A2(n19), .ZN(n63) );
  nr02d0 U49 ( .A1(n24), .A2(n20), .ZN(n64) );
  nr02d0 U50 ( .A1(n25), .A2(n20), .ZN(n65) );
  nr02d0 U51 ( .A1(n26), .A2(n20), .ZN(n66) );
  nr02d0 U52 ( .A1(n27), .A2(n20), .ZN(n67) );
  nr02d0 U53 ( .A1(n28), .A2(n20), .ZN(n68) );
  nr02d0 U54 ( .A1(n29), .A2(n20), .ZN(n69) );
  nr02d0 U55 ( .A1(n30), .A2(n20), .ZN(n70) );
  nr02d0 U56 ( .A1(n31), .A2(n20), .ZN(n71) );
  nr02d0 U57 ( .A1(n24), .A2(n21), .ZN(n72) );
  nr02d0 U58 ( .A1(n25), .A2(n21), .ZN(n73) );
  nr02d0 U59 ( .A1(n26), .A2(n21), .ZN(n74) );
  nr02d0 U60 ( .A1(n27), .A2(n21), .ZN(n75) );
  nr02d0 U61 ( .A1(n28), .A2(n21), .ZN(n76) );
  nr02d0 U62 ( .A1(n29), .A2(n21), .ZN(n77) );
  nr02d0 U63 ( .A1(n30), .A2(n21), .ZN(n78) );
  nr02d0 U64 ( .A1(n31), .A2(n21), .ZN(n79) );
  nr02d0 U65 ( .A1(n24), .A2(n22), .ZN(n80) );
  nr02d0 U66 ( .A1(n25), .A2(n22), .ZN(n81) );
  nr02d0 U67 ( .A1(n26), .A2(n22), .ZN(n82) );
  nr02d0 U68 ( .A1(n27), .A2(n22), .ZN(n83) );
  nr02d0 U69 ( .A1(n28), .A2(n22), .ZN(n84) );
  nr02d0 U70 ( .A1(n29), .A2(n22), .ZN(n85) );
  nr02d0 U71 ( .A1(n30), .A2(n22), .ZN(n86) );
  nr02d0 U72 ( .A1(n31), .A2(n22), .ZN(n87) );
  nr02d0 U73 ( .A1(n24), .A2(n23), .ZN(n88) );
  nr02d0 U74 ( .A1(n25), .A2(n23), .ZN(n89) );
  nr02d0 U75 ( .A1(n26), .A2(n23), .ZN(n90) );
  nr02d0 U76 ( .A1(n27), .A2(n23), .ZN(n91) );
  nr02d0 U77 ( .A1(n28), .A2(n23), .ZN(n92) );
  nr02d0 U78 ( .A1(n29), .A2(n23), .ZN(n93) );
  nr02d0 U79 ( .A1(n30), .A2(n23), .ZN(n94) );
  nr02d0 U80 ( .A1(n31), .A2(n23), .ZN(n95) );
  ah01d0 U81 ( .A(n34), .B(n41), .CO(n97), .S(n96) );
  ah01d0 U82 ( .A(n49), .B(n56), .CO(n99), .S(n98) );
  ad01d0 U83 ( .A(n35), .B(n42), .CI(n97), .CO(n101), .S(n100) );
  ah01d0 U84 ( .A(n57), .B(n64), .CO(n103), .S(n102) );
  ad01d0 U85 ( .A(n36), .B(n50), .CI(n43), .CO(n105), .S(n104) );
  ad01d0 U86 ( .A(n99), .B(n102), .CI(n104), .CO(n107), .S(n106) );
  ah01d0 U87 ( .A(n65), .B(n72), .CO(n109), .S(n108) );
  ad01d0 U88 ( .A(n37), .B(n58), .CI(n51), .CO(n111), .S(n110) );
  ad01d0 U89 ( .A(n44), .B(n103), .CI(n108), .CO(n113), .S(n112) );
  ad01d0 U90 ( .A(n105), .B(n110), .CI(n112), .CO(n115), .S(n114) );
  ah01d0 U91 ( .A(n73), .B(n80), .CO(n117), .S(n116) );
  ad01d0 U92 ( .A(n38), .B(n66), .CI(n45), .CO(n119), .S(n118) );
  ad01d0 U93 ( .A(n52), .B(n59), .CI(n109), .CO(n121), .S(n120) );
  ad01d0 U94 ( .A(n116), .B(n111), .CI(n118), .CO(n123), .S(n122) );
  ad01d0 U95 ( .A(n113), .B(n120), .CI(n122), .CO(n125), .S(n124) );
  ah01d0 U96 ( .A(n81), .B(n88), .CO(n127), .S(n126) );
  ad01d0 U97 ( .A(n39), .B(n74), .CI(n46), .CO(n129), .S(n128) );
  ad01d0 U98 ( .A(n53), .B(n67), .CI(n60), .CO(n131), .S(n130) );
  ad01d0 U99 ( .A(n117), .B(n126), .CI(n119), .CO(n133), .S(n132) );
  ad01d0 U100 ( .A(n130), .B(n128), .CI(n121), .CO(n135), .S(n134) );
  ad01d0 U101 ( .A(n132), .B(n123), .CI(n134), .CO(n137), .S(n136) );
  ah01d0 U102 ( .A(n82), .B(n89), .CO(n139), .S(n138) );
  ad01d0 U103 ( .A(n68), .B(n75), .CI(n47), .CO(n141), .S(n140) );
  ad01d0 U104 ( .A(n54), .B(n61), .CI(n127), .CO(n143), .S(n142) );
  ad01d0 U105 ( .A(n138), .B(n129), .CI(n131), .CO(n145), .S(n144) );
  ad01d0 U106 ( .A(n140), .B(n142), .CI(n133), .CO(n147), .S(n146) );
  ad01d0 U107 ( .A(n144), .B(n135), .CI(n146), .CO(n149), .S(n148) );
  ad01d0 U108 ( .A(n55), .B(n90), .CI(n83), .CO(n151), .S(n150) );
  ad01d0 U109 ( .A(n76), .B(n69), .CI(n62), .CO(n153), .S(n152) );
  ad01d0 U110 ( .A(n139), .B(n141), .CI(n152), .CO(n155), .S(n154) );
  ad01d0 U111 ( .A(n150), .B(n143), .CI(n145), .CO(n157), .S(n156) );
  ad01d0 U112 ( .A(n154), .B(n147), .CI(n156), .CO(n159), .S(n158) );
  ad01d0 U113 ( .A(n63), .B(n91), .CI(n84), .CO(n161), .S(n160) );
  ad01d0 U114 ( .A(n70), .B(n77), .CI(n151), .CO(n163), .S(n162) );
  ad01d0 U115 ( .A(n153), .B(n160), .CI(n162), .CO(n165), .S(n164) );
  ad01d0 U116 ( .A(n155), .B(n157), .CI(n164), .CO(n167), .S(n166) );
  ad01d0 U117 ( .A(n71), .B(n92), .CI(n85), .CO(n169), .S(n168) );
  ad01d0 U118 ( .A(n78), .B(n161), .CI(n168), .CO(n171), .S(n170) );
  ad01d0 U119 ( .A(n163), .B(n170), .CI(n165), .CO(n173), .S(n172) );
  ad01d0 U120 ( .A(n79), .B(n93), .CI(n86), .CO(n175), .S(n174) );
  ad01d0 U121 ( .A(n169), .B(n174), .CI(n171), .CO(n177), .S(n176) );
  ad01d0 U122 ( .A(n87), .B(n94), .CI(n175), .CO(n179), .S(n178) );
  ah01d0 U123 ( .A(n40), .B(n33), .CO(n180), .S(product[1]) );
  ad01d0 U124 ( .A(n48), .B(n180), .CI(n96), .CO(n181), .S(product[2]) );
  ad01d0 U125 ( .A(n98), .B(n181), .CI(n100), .CO(n182), .S(product[3]) );
  ad01d0 U126 ( .A(n101), .B(n106), .CI(n182), .CO(n183), .S(product[4]) );
  ad01d0 U127 ( .A(n107), .B(n114), .CI(n183), .CO(n184), .S(product[5]) );
  ad01d0 U128 ( .A(n115), .B(n124), .CI(n184), .CO(n185), .S(product[6]) );
  ad01d0 U129 ( .A(n125), .B(n136), .CI(n185), .CO(n186), .S(product[7]) );
  ad01d0 U130 ( .A(n137), .B(n148), .CI(n186), .CO(n187), .S(product[8]) );
  ad01d0 U131 ( .A(n149), .B(n158), .CI(n187), .CO(n188), .S(product[9]) );
  ad01d0 U132 ( .A(n159), .B(n166), .CI(n188), .CO(n189), .S(product[10]) );
  ad01d0 U133 ( .A(n167), .B(n172), .CI(n189), .CO(n190), .S(product[11]) );
  ad01d0 U134 ( .A(n176), .B(n173), .CI(n190), .CO(n191), .S(product[12]) );
  ad01d0 U135 ( .A(n178), .B(n177), .CI(n191), .CO(n192), .S(product[13]) );
  ad01d0 U136 ( .A(n95), .B(n179), .CI(n192), .CO(product[15]), .S(product[14]) );
  inv0d1 U140 ( .I(a[4]), .ZN(n20) );
  inv0d1 U141 ( .I(a[3]), .ZN(n19) );
  inv0d1 U142 ( .I(a[0]), .ZN(n16) );
  inv0d1 U143 ( .I(a[2]), .ZN(n18) );
  inv0d1 U144 ( .I(a[1]), .ZN(n17) );
  inv0d1 U145 ( .I(a[5]), .ZN(n21) );
  inv0d1 U146 ( .I(a[6]), .ZN(n22) );
  inv0d1 U147 ( .I(a[7]), .ZN(n23) );
  inv0d1 U148 ( .I(b[1]), .ZN(n25) );
  inv0d1 U149 ( .I(b[0]), .ZN(n24) );
  inv0d1 U150 ( .I(b[2]), .ZN(n26) );
  inv0d1 U151 ( .I(b[3]), .ZN(n27) );
  inv0d1 U152 ( .I(b[4]), .ZN(n28) );
  inv0d1 U153 ( .I(b[5]), .ZN(n29) );
  inv0d1 U154 ( .I(b[6]), .ZN(n30) );
  inv0d1 U155 ( .I(b[7]), .ZN(n31) );
endmodule


module SDRAM_FIFO_1 ( fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, 
        fifo_push_req_n, fifo_pop_req_n, fifo_data_in, push_empty_fifo, 
        push_ae_fifo, push_hf_fifo, push_af_fifo, push_full_fifo, 
        push_error_fifo, pop_empty_fifo, pop_ae_fifo, pop_hf_fifo, pop_af_fifo, 
        pop_full_fifo, pop_error_fifo, data_out_fifo, test_se, test_si1, 
        test_si2, test_so1, test_so2 );
  input [31:0] fifo_data_in;
  output [31:0] data_out_fifo;
  input fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, fifo_push_req_n,
         fifo_pop_req_n, test_se, test_si1, test_si2;
  output push_empty_fifo, push_ae_fifo, push_hf_fifo, push_af_fifo,
         push_full_fifo, push_error_fifo, pop_empty_fifo, pop_ae_fifo,
         pop_hf_fifo, pop_af_fifo, pop_full_fifo, pop_error_fifo, test_so1,
         test_so2;
  wire   we_n, wr_addr_2_, wr_addr_1_, wr_addr_0_, rd_addr_2_, rd_addr_1_,
         rd_addr_0_, reg_array_0__31_, reg_array_0__30_, reg_array_0__29_,
         reg_array_0__28_, reg_array_0__27_, reg_array_0__26_,
         reg_array_0__25_, reg_array_0__24_, reg_array_0__23_,
         reg_array_0__22_, reg_array_0__21_, reg_array_0__20_,
         reg_array_0__19_, reg_array_0__18_, reg_array_0__17_,
         reg_array_0__16_, reg_array_0__15_, reg_array_0__14_,
         reg_array_0__13_, reg_array_0__12_, reg_array_0__11_,
         reg_array_0__10_, reg_array_0__9_, reg_array_0__8_, reg_array_0__7_,
         reg_array_0__6_, reg_array_0__5_, reg_array_0__4_, reg_array_0__3_,
         reg_array_0__2_, reg_array_0__1_, reg_array_0__0_, reg_array_1__31_,
         reg_array_1__30_, reg_array_1__29_, reg_array_1__28_,
         reg_array_1__27_, reg_array_1__26_, reg_array_1__25_,
         reg_array_1__24_, reg_array_1__23_, reg_array_1__22_,
         reg_array_1__21_, reg_array_1__20_, reg_array_1__19_,
         reg_array_1__18_, reg_array_1__17_, reg_array_1__16_,
         reg_array_1__15_, reg_array_1__14_, reg_array_1__13_,
         reg_array_1__12_, reg_array_1__11_, reg_array_1__10_, reg_array_1__9_,
         reg_array_1__8_, reg_array_1__7_, reg_array_1__6_, reg_array_1__5_,
         reg_array_1__4_, reg_array_1__3_, reg_array_1__2_, reg_array_1__1_,
         reg_array_1__0_, reg_array_2__31_, reg_array_2__30_, reg_array_2__29_,
         reg_array_2__28_, reg_array_2__27_, reg_array_2__26_,
         reg_array_2__25_, reg_array_2__24_, reg_array_2__23_,
         reg_array_2__22_, reg_array_2__21_, reg_array_2__20_,
         reg_array_2__19_, reg_array_2__18_, reg_array_2__17_,
         reg_array_2__16_, reg_array_2__15_, reg_array_2__14_,
         reg_array_2__13_, reg_array_2__12_, reg_array_2__11_,
         reg_array_2__10_, reg_array_2__9_, reg_array_2__8_, reg_array_2__7_,
         reg_array_2__6_, reg_array_2__5_, reg_array_2__4_, reg_array_2__3_,
         reg_array_2__2_, reg_array_2__1_, reg_array_2__0_, reg_array_3__31_,
         reg_array_3__30_, reg_array_3__29_, reg_array_3__28_,
         reg_array_3__27_, reg_array_3__26_, reg_array_3__25_,
         reg_array_3__24_, reg_array_3__23_, reg_array_3__22_,
         reg_array_3__21_, reg_array_3__20_, reg_array_3__19_,
         reg_array_3__18_, reg_array_3__17_, reg_array_3__16_,
         reg_array_3__15_, reg_array_3__14_, reg_array_3__13_,
         reg_array_3__12_, reg_array_3__11_, reg_array_3__10_, reg_array_3__9_,
         reg_array_3__8_, reg_array_3__7_, reg_array_3__6_, reg_array_3__5_,
         reg_array_3__4_, reg_array_3__3_, reg_array_3__2_, reg_array_3__1_,
         reg_array_3__0_, reg_array_4__31_, reg_array_4__30_, reg_array_4__29_,
         reg_array_4__28_, reg_array_4__27_, reg_array_4__26_,
         reg_array_4__25_, reg_array_4__24_, reg_array_4__23_,
         reg_array_4__22_, reg_array_4__21_, reg_array_4__20_,
         reg_array_4__19_, reg_array_4__18_, reg_array_4__17_,
         reg_array_4__16_, reg_array_4__15_, reg_array_4__14_,
         reg_array_4__13_, reg_array_4__12_, reg_array_4__11_,
         reg_array_4__10_, reg_array_4__9_, reg_array_4__8_, reg_array_4__7_,
         reg_array_4__6_, reg_array_4__5_, reg_array_4__4_, reg_array_4__3_,
         reg_array_4__2_, reg_array_4__1_, reg_array_4__0_, reg_array_5__31_,
         reg_array_5__30_, reg_array_5__29_, reg_array_5__28_,
         reg_array_5__27_, reg_array_5__26_, reg_array_5__25_,
         reg_array_5__24_, reg_array_5__23_, reg_array_5__22_,
         reg_array_5__21_, reg_array_5__20_, reg_array_5__19_,
         reg_array_5__18_, reg_array_5__17_, reg_array_5__16_,
         reg_array_5__15_, reg_array_5__14_, reg_array_5__13_,
         reg_array_5__12_, reg_array_5__11_, reg_array_5__10_, reg_array_5__9_,
         reg_array_5__8_, reg_array_5__7_, reg_array_5__6_, reg_array_5__5_,
         reg_array_5__4_, reg_array_5__3_, reg_array_5__2_, reg_array_5__1_,
         reg_array_5__0_, reg_array_6__31_, reg_array_6__30_, reg_array_6__29_,
         reg_array_6__28_, reg_array_6__27_, reg_array_6__26_,
         reg_array_6__25_, reg_array_6__24_, reg_array_6__23_,
         reg_array_6__22_, reg_array_6__21_, reg_array_6__20_,
         reg_array_6__19_, reg_array_6__18_, reg_array_6__17_,
         reg_array_6__16_, reg_array_6__15_, reg_array_6__14_,
         reg_array_6__13_, reg_array_6__12_, reg_array_6__11_,
         reg_array_6__10_, reg_array_6__9_, reg_array_6__8_, reg_array_6__7_,
         reg_array_6__6_, reg_array_6__5_, reg_array_6__4_, reg_array_6__3_,
         reg_array_6__2_, reg_array_6__1_, reg_array_6__0_, reg_array_7__30_,
         reg_array_7__29_, reg_array_7__28_, reg_array_7__27_,
         reg_array_7__26_, reg_array_7__25_, reg_array_7__24_,
         reg_array_7__23_, reg_array_7__22_, reg_array_7__21_,
         reg_array_7__20_, reg_array_7__19_, reg_array_7__18_,
         reg_array_7__17_, reg_array_7__16_, reg_array_7__15_,
         reg_array_7__14_, reg_array_7__13_, reg_array_7__12_,
         reg_array_7__11_, reg_array_7__10_, reg_array_7__9_, reg_array_7__8_,
         reg_array_7__7_, reg_array_7__6_, reg_array_7__5_, reg_array_7__4_,
         reg_array_7__3_, reg_array_7__2_, reg_array_7__1_, reg_array_7__0_,
         N729, N731, N733, N735, N737, N739, N741, N743, N745, N747, N749,
         N751, N753, N755, N757, N759, N761, N763, N765, N767, N769, N771,
         N773, N775, N777, N779, N781, N783, N785, N787, N789, N791, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838,
         data_out_sync_31_, data_out_sync_30_, data_out_sync_29_,
         data_out_sync_28_, data_out_sync_27_, data_out_sync_26_,
         data_out_sync_25_, data_out_sync_24_, data_out_sync_23_,
         data_out_sync_22_, data_out_sync_21_, data_out_sync_20_,
         data_out_sync_19_, data_out_sync_18_, data_out_sync_17_,
         data_out_sync_16_, data_out_sync_15_, data_out_sync_14_,
         data_out_sync_13_, data_out_sync_12_, data_out_sync_11_,
         data_out_sync_10_, data_out_sync_9_, data_out_sync_8_,
         data_out_sync_7_, data_out_sync_6_, data_out_sync_5_,
         data_out_sync_4_, data_out_sync_3_, data_out_sync_2_,
         data_out_sync_1_, data_out_sync_0_, n1, n97, n130, n163, n196, n229,
         n262, n295, n328, n404, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n869, n872, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16;

  an03d1 U363 ( .A1(n475), .A2(n474), .A3(rd_addr_2_), .Z(n542) );
  an03d1 U364 ( .A1(rd_addr_0_), .A2(n474), .A3(rd_addr_2_), .Z(n543) );
  an03d1 U365 ( .A1(rd_addr_1_), .A2(n475), .A3(rd_addr_2_), .Z(n544) );
  an03d1 U366 ( .A1(rd_addr_1_), .A2(rd_addr_0_), .A3(rd_addr_2_), .Z(n545) );
  an02d1 U379 ( .A1(fifo_rst_n), .A2(fifo_data_in[31]), .Z(N791) );
  an02d1 U380 ( .A1(fifo_data_in[30]), .A2(fifo_rst_n), .Z(N789) );
  an02d1 U381 ( .A1(fifo_data_in[29]), .A2(fifo_rst_n), .Z(N787) );
  an02d1 U382 ( .A1(fifo_data_in[28]), .A2(fifo_rst_n), .Z(N785) );
  an02d1 U383 ( .A1(fifo_data_in[27]), .A2(fifo_rst_n), .Z(N783) );
  an02d1 U384 ( .A1(fifo_data_in[26]), .A2(fifo_rst_n), .Z(N781) );
  an02d1 U385 ( .A1(fifo_data_in[25]), .A2(fifo_rst_n), .Z(N779) );
  an02d1 U386 ( .A1(fifo_data_in[24]), .A2(fifo_rst_n), .Z(N777) );
  an02d1 U387 ( .A1(fifo_data_in[23]), .A2(fifo_rst_n), .Z(N775) );
  an02d1 U388 ( .A1(fifo_data_in[22]), .A2(fifo_rst_n), .Z(N773) );
  an02d1 U389 ( .A1(fifo_data_in[21]), .A2(fifo_rst_n), .Z(N771) );
  an02d1 U390 ( .A1(fifo_data_in[20]), .A2(fifo_rst_n), .Z(N769) );
  an02d1 U391 ( .A1(fifo_data_in[19]), .A2(fifo_rst_n), .Z(N767) );
  an02d1 U392 ( .A1(fifo_data_in[18]), .A2(fifo_rst_n), .Z(N765) );
  an02d1 U393 ( .A1(fifo_data_in[17]), .A2(fifo_rst_n), .Z(N763) );
  an02d1 U394 ( .A1(fifo_data_in[16]), .A2(fifo_rst_n), .Z(N761) );
  an02d1 U395 ( .A1(fifo_data_in[15]), .A2(fifo_rst_n), .Z(N759) );
  an02d1 U396 ( .A1(fifo_data_in[14]), .A2(fifo_rst_n), .Z(N757) );
  an02d1 U397 ( .A1(fifo_data_in[13]), .A2(fifo_rst_n), .Z(N755) );
  an02d1 U398 ( .A1(fifo_data_in[12]), .A2(fifo_rst_n), .Z(N753) );
  an02d1 U399 ( .A1(fifo_data_in[11]), .A2(fifo_rst_n), .Z(N751) );
  an02d1 U400 ( .A1(fifo_data_in[10]), .A2(fifo_rst_n), .Z(N749) );
  an02d1 U401 ( .A1(fifo_data_in[9]), .A2(fifo_rst_n), .Z(N747) );
  an02d1 U402 ( .A1(fifo_data_in[8]), .A2(fifo_rst_n), .Z(N745) );
  an02d1 U403 ( .A1(fifo_data_in[7]), .A2(fifo_rst_n), .Z(N743) );
  an02d1 U404 ( .A1(fifo_data_in[6]), .A2(fifo_rst_n), .Z(N741) );
  an02d1 U405 ( .A1(fifo_data_in[5]), .A2(fifo_rst_n), .Z(N739) );
  an02d1 U406 ( .A1(fifo_data_in[4]), .A2(fifo_rst_n), .Z(N737) );
  an02d1 U407 ( .A1(fifo_data_in[3]), .A2(fifo_rst_n), .Z(N735) );
  an02d1 U408 ( .A1(fifo_data_in[2]), .A2(fifo_rst_n), .Z(N733) );
  an02d1 U409 ( .A1(fifo_data_in[1]), .A2(fifo_rst_n), .Z(N731) );
  an02d1 U410 ( .A1(fifo_data_in[0]), .A2(fifo_rst_n), .Z(N729) );
  aoi2222d1 U413 ( .A1(reg_array_7__0_), .A2(n438), .B1(reg_array_6__0_), .B2(
        n435), .C1(reg_array_5__0_), .C2(n432), .D1(reg_array_4__0_), .D2(n429), .ZN(n546) );
  aoi2222d1 U414 ( .A1(reg_array_3__0_), .A2(n426), .B1(reg_array_2__0_), .B2(
        n423), .C1(reg_array_1__0_), .C2(n420), .D1(reg_array_0__0_), .D2(n417), .ZN(n547) );
  aoi2222d1 U415 ( .A1(reg_array_7__1_), .A2(n438), .B1(reg_array_6__1_), .B2(
        n435), .C1(reg_array_5__1_), .C2(n432), .D1(reg_array_4__1_), .D2(n429), .ZN(n536) );
  aoi2222d1 U416 ( .A1(reg_array_3__1_), .A2(n426), .B1(reg_array_2__1_), .B2(
        n423), .C1(reg_array_1__1_), .C2(n420), .D1(reg_array_0__1_), .D2(n417), .ZN(n537) );
  aoi2222d1 U417 ( .A1(reg_array_7__2_), .A2(n438), .B1(reg_array_6__2_), .B2(
        n435), .C1(reg_array_5__2_), .C2(n432), .D1(reg_array_4__2_), .D2(n429), .ZN(n534) );
  aoi2222d1 U418 ( .A1(reg_array_3__2_), .A2(n426), .B1(reg_array_2__2_), .B2(
        n423), .C1(reg_array_1__2_), .C2(n420), .D1(reg_array_0__2_), .D2(n417), .ZN(n535) );
  aoi2222d1 U419 ( .A1(reg_array_7__3_), .A2(n438), .B1(reg_array_6__3_), .B2(
        n435), .C1(reg_array_5__3_), .C2(n432), .D1(reg_array_4__3_), .D2(n429), .ZN(n532) );
  aoi2222d1 U420 ( .A1(reg_array_3__3_), .A2(n426), .B1(reg_array_2__3_), .B2(
        n423), .C1(reg_array_1__3_), .C2(n420), .D1(reg_array_0__3_), .D2(n417), .ZN(n533) );
  aoi2222d1 U421 ( .A1(reg_array_7__4_), .A2(n438), .B1(reg_array_6__4_), .B2(
        n435), .C1(reg_array_5__4_), .C2(n432), .D1(reg_array_4__4_), .D2(n429), .ZN(n530) );
  aoi2222d1 U422 ( .A1(reg_array_3__4_), .A2(n426), .B1(reg_array_2__4_), .B2(
        n423), .C1(reg_array_1__4_), .C2(n420), .D1(reg_array_0__4_), .D2(n417), .ZN(n531) );
  aoi2222d1 U423 ( .A1(reg_array_7__5_), .A2(n438), .B1(reg_array_6__5_), .B2(
        n435), .C1(reg_array_5__5_), .C2(n432), .D1(reg_array_4__5_), .D2(n429), .ZN(n528) );
  aoi2222d1 U424 ( .A1(reg_array_3__5_), .A2(n426), .B1(reg_array_2__5_), .B2(
        n423), .C1(reg_array_1__5_), .C2(n420), .D1(reg_array_0__5_), .D2(n417), .ZN(n529) );
  aoi2222d1 U425 ( .A1(reg_array_7__6_), .A2(n438), .B1(reg_array_6__6_), .B2(
        n435), .C1(reg_array_5__6_), .C2(n432), .D1(reg_array_4__6_), .D2(n429), .ZN(n526) );
  aoi2222d1 U426 ( .A1(reg_array_3__6_), .A2(n426), .B1(reg_array_2__6_), .B2(
        n423), .C1(reg_array_1__6_), .C2(n420), .D1(reg_array_0__6_), .D2(n417), .ZN(n527) );
  aoi2222d1 U427 ( .A1(reg_array_7__7_), .A2(n438), .B1(reg_array_6__7_), .B2(
        n435), .C1(reg_array_5__7_), .C2(n432), .D1(reg_array_4__7_), .D2(n429), .ZN(n524) );
  aoi2222d1 U428 ( .A1(reg_array_3__7_), .A2(n426), .B1(reg_array_2__7_), .B2(
        n423), .C1(reg_array_1__7_), .C2(n420), .D1(reg_array_0__7_), .D2(n417), .ZN(n525) );
  aoi2222d1 U429 ( .A1(reg_array_7__8_), .A2(n438), .B1(reg_array_6__8_), .B2(
        n435), .C1(reg_array_5__8_), .C2(n432), .D1(reg_array_4__8_), .D2(n429), .ZN(n522) );
  aoi2222d1 U430 ( .A1(reg_array_3__8_), .A2(n426), .B1(reg_array_2__8_), .B2(
        n423), .C1(reg_array_1__8_), .C2(n420), .D1(reg_array_0__8_), .D2(n417), .ZN(n523) );
  aoi2222d1 U431 ( .A1(reg_array_7__9_), .A2(n438), .B1(reg_array_6__9_), .B2(
        n435), .C1(reg_array_5__9_), .C2(n432), .D1(reg_array_4__9_), .D2(n429), .ZN(n520) );
  aoi2222d1 U432 ( .A1(reg_array_3__9_), .A2(n426), .B1(reg_array_2__9_), .B2(
        n423), .C1(reg_array_1__9_), .C2(n420), .D1(reg_array_0__9_), .D2(n417), .ZN(n521) );
  aoi2222d1 U433 ( .A1(reg_array_7__10_), .A2(n437), .B1(reg_array_6__10_), 
        .B2(n434), .C1(reg_array_5__10_), .C2(n431), .D1(reg_array_4__10_), 
        .D2(n428), .ZN(n518) );
  aoi2222d1 U434 ( .A1(reg_array_3__10_), .A2(n425), .B1(reg_array_2__10_), 
        .B2(n422), .C1(reg_array_1__10_), .C2(n419), .D1(reg_array_0__10_), 
        .D2(n416), .ZN(n519) );
  aoi2222d1 U435 ( .A1(reg_array_7__11_), .A2(n437), .B1(reg_array_6__11_), 
        .B2(n434), .C1(reg_array_5__11_), .C2(n431), .D1(reg_array_4__11_), 
        .D2(n428), .ZN(n516) );
  aoi2222d1 U436 ( .A1(reg_array_3__11_), .A2(n425), .B1(reg_array_2__11_), 
        .B2(n422), .C1(reg_array_1__11_), .C2(n419), .D1(reg_array_0__11_), 
        .D2(n416), .ZN(n517) );
  aoi2222d1 U437 ( .A1(reg_array_7__12_), .A2(n437), .B1(reg_array_6__12_), 
        .B2(n434), .C1(reg_array_5__12_), .C2(n431), .D1(reg_array_4__12_), 
        .D2(n428), .ZN(n514) );
  aoi2222d1 U438 ( .A1(reg_array_3__12_), .A2(n425), .B1(reg_array_2__12_), 
        .B2(n422), .C1(reg_array_1__12_), .C2(n419), .D1(reg_array_0__12_), 
        .D2(n416), .ZN(n515) );
  aoi2222d1 U439 ( .A1(reg_array_7__13_), .A2(n437), .B1(reg_array_6__13_), 
        .B2(n434), .C1(reg_array_5__13_), .C2(n431), .D1(reg_array_4__13_), 
        .D2(n428), .ZN(n512) );
  aoi2222d1 U440 ( .A1(reg_array_3__13_), .A2(n425), .B1(reg_array_2__13_), 
        .B2(n422), .C1(reg_array_1__13_), .C2(n419), .D1(reg_array_0__13_), 
        .D2(n416), .ZN(n513) );
  aoi2222d1 U441 ( .A1(reg_array_7__14_), .A2(n437), .B1(reg_array_6__14_), 
        .B2(n434), .C1(reg_array_5__14_), .C2(n431), .D1(reg_array_4__14_), 
        .D2(n428), .ZN(n510) );
  aoi2222d1 U442 ( .A1(reg_array_3__14_), .A2(n425), .B1(reg_array_2__14_), 
        .B2(n422), .C1(reg_array_1__14_), .C2(n419), .D1(reg_array_0__14_), 
        .D2(n416), .ZN(n511) );
  aoi2222d1 U443 ( .A1(reg_array_7__15_), .A2(n437), .B1(reg_array_6__15_), 
        .B2(n434), .C1(reg_array_5__15_), .C2(n431), .D1(reg_array_4__15_), 
        .D2(n428), .ZN(n508) );
  aoi2222d1 U444 ( .A1(reg_array_3__15_), .A2(n425), .B1(reg_array_2__15_), 
        .B2(n422), .C1(reg_array_1__15_), .C2(n419), .D1(reg_array_0__15_), 
        .D2(n416), .ZN(n509) );
  aoi2222d1 U445 ( .A1(reg_array_7__16_), .A2(n437), .B1(reg_array_6__16_), 
        .B2(n434), .C1(reg_array_5__16_), .C2(n431), .D1(reg_array_4__16_), 
        .D2(n428), .ZN(n506) );
  aoi2222d1 U446 ( .A1(reg_array_3__16_), .A2(n425), .B1(reg_array_2__16_), 
        .B2(n422), .C1(reg_array_1__16_), .C2(n419), .D1(reg_array_0__16_), 
        .D2(n416), .ZN(n507) );
  aoi2222d1 U447 ( .A1(reg_array_7__17_), .A2(n437), .B1(reg_array_6__17_), 
        .B2(n434), .C1(reg_array_5__17_), .C2(n431), .D1(reg_array_4__17_), 
        .D2(n428), .ZN(n504) );
  aoi2222d1 U448 ( .A1(reg_array_3__17_), .A2(n425), .B1(reg_array_2__17_), 
        .B2(n422), .C1(reg_array_1__17_), .C2(n419), .D1(reg_array_0__17_), 
        .D2(n416), .ZN(n505) );
  aoi2222d1 U449 ( .A1(reg_array_7__18_), .A2(n437), .B1(reg_array_6__18_), 
        .B2(n434), .C1(reg_array_5__18_), .C2(n431), .D1(reg_array_4__18_), 
        .D2(n428), .ZN(n502) );
  aoi2222d1 U450 ( .A1(reg_array_3__18_), .A2(n425), .B1(reg_array_2__18_), 
        .B2(n422), .C1(reg_array_1__18_), .C2(n419), .D1(reg_array_0__18_), 
        .D2(n416), .ZN(n503) );
  aoi2222d1 U451 ( .A1(reg_array_7__19_), .A2(n437), .B1(reg_array_6__19_), 
        .B2(n434), .C1(reg_array_5__19_), .C2(n431), .D1(reg_array_4__19_), 
        .D2(n428), .ZN(n500) );
  aoi2222d1 U452 ( .A1(reg_array_3__19_), .A2(n425), .B1(reg_array_2__19_), 
        .B2(n422), .C1(reg_array_1__19_), .C2(n419), .D1(reg_array_0__19_), 
        .D2(n416), .ZN(n501) );
  aoi2222d1 U453 ( .A1(reg_array_7__20_), .A2(n437), .B1(reg_array_6__20_), 
        .B2(n434), .C1(reg_array_5__20_), .C2(n431), .D1(reg_array_4__20_), 
        .D2(n428), .ZN(n498) );
  aoi2222d1 U454 ( .A1(reg_array_3__20_), .A2(n425), .B1(reg_array_2__20_), 
        .B2(n422), .C1(reg_array_1__20_), .C2(n419), .D1(reg_array_0__20_), 
        .D2(n416), .ZN(n499) );
  aoi2222d1 U455 ( .A1(reg_array_7__21_), .A2(n436), .B1(reg_array_6__21_), 
        .B2(n433), .C1(reg_array_5__21_), .C2(n430), .D1(reg_array_4__21_), 
        .D2(n427), .ZN(n496) );
  aoi2222d1 U456 ( .A1(reg_array_3__21_), .A2(n424), .B1(reg_array_2__21_), 
        .B2(n421), .C1(reg_array_1__21_), .C2(n418), .D1(reg_array_0__21_), 
        .D2(n404), .ZN(n497) );
  aoi2222d1 U457 ( .A1(reg_array_7__22_), .A2(n436), .B1(reg_array_6__22_), 
        .B2(n433), .C1(reg_array_5__22_), .C2(n430), .D1(reg_array_4__22_), 
        .D2(n427), .ZN(n494) );
  aoi2222d1 U458 ( .A1(reg_array_3__22_), .A2(n424), .B1(reg_array_2__22_), 
        .B2(n421), .C1(reg_array_1__22_), .C2(n418), .D1(reg_array_0__22_), 
        .D2(n404), .ZN(n495) );
  aoi2222d1 U459 ( .A1(reg_array_7__23_), .A2(n436), .B1(reg_array_6__23_), 
        .B2(n433), .C1(reg_array_5__23_), .C2(n430), .D1(reg_array_4__23_), 
        .D2(n427), .ZN(n492) );
  aoi2222d1 U460 ( .A1(reg_array_3__23_), .A2(n424), .B1(reg_array_2__23_), 
        .B2(n421), .C1(reg_array_1__23_), .C2(n418), .D1(reg_array_0__23_), 
        .D2(n404), .ZN(n493) );
  aoi2222d1 U461 ( .A1(reg_array_7__24_), .A2(n436), .B1(reg_array_6__24_), 
        .B2(n433), .C1(reg_array_5__24_), .C2(n430), .D1(reg_array_4__24_), 
        .D2(n427), .ZN(n490) );
  aoi2222d1 U462 ( .A1(reg_array_3__24_), .A2(n424), .B1(reg_array_2__24_), 
        .B2(n421), .C1(reg_array_1__24_), .C2(n418), .D1(reg_array_0__24_), 
        .D2(n404), .ZN(n491) );
  aoi2222d1 U463 ( .A1(reg_array_7__25_), .A2(n436), .B1(reg_array_6__25_), 
        .B2(n433), .C1(reg_array_5__25_), .C2(n430), .D1(reg_array_4__25_), 
        .D2(n427), .ZN(n488) );
  aoi2222d1 U464 ( .A1(reg_array_3__25_), .A2(n424), .B1(reg_array_2__25_), 
        .B2(n421), .C1(reg_array_1__25_), .C2(n418), .D1(reg_array_0__25_), 
        .D2(n404), .ZN(n489) );
  aoi2222d1 U465 ( .A1(reg_array_7__26_), .A2(n436), .B1(reg_array_6__26_), 
        .B2(n433), .C1(reg_array_5__26_), .C2(n430), .D1(reg_array_4__26_), 
        .D2(n427), .ZN(n486) );
  aoi2222d1 U466 ( .A1(reg_array_3__26_), .A2(n424), .B1(reg_array_2__26_), 
        .B2(n421), .C1(reg_array_1__26_), .C2(n418), .D1(reg_array_0__26_), 
        .D2(n404), .ZN(n487) );
  aoi2222d1 U467 ( .A1(reg_array_7__27_), .A2(n436), .B1(reg_array_6__27_), 
        .B2(n433), .C1(reg_array_5__27_), .C2(n430), .D1(reg_array_4__27_), 
        .D2(n427), .ZN(n484) );
  aoi2222d1 U468 ( .A1(reg_array_3__27_), .A2(n424), .B1(reg_array_2__27_), 
        .B2(n421), .C1(reg_array_1__27_), .C2(n418), .D1(reg_array_0__27_), 
        .D2(n404), .ZN(n485) );
  aoi2222d1 U469 ( .A1(reg_array_7__28_), .A2(n436), .B1(reg_array_6__28_), 
        .B2(n433), .C1(reg_array_5__28_), .C2(n430), .D1(reg_array_4__28_), 
        .D2(n427), .ZN(n482) );
  aoi2222d1 U470 ( .A1(reg_array_3__28_), .A2(n424), .B1(reg_array_2__28_), 
        .B2(n421), .C1(reg_array_1__28_), .C2(n418), .D1(reg_array_0__28_), 
        .D2(n404), .ZN(n483) );
  aoi2222d1 U471 ( .A1(reg_array_7__29_), .A2(n436), .B1(reg_array_6__29_), 
        .B2(n433), .C1(reg_array_5__29_), .C2(n430), .D1(reg_array_4__29_), 
        .D2(n427), .ZN(n480) );
  aoi2222d1 U472 ( .A1(reg_array_3__29_), .A2(n424), .B1(reg_array_2__29_), 
        .B2(n421), .C1(reg_array_1__29_), .C2(n418), .D1(reg_array_0__29_), 
        .D2(n404), .ZN(n481) );
  aoi2222d1 U473 ( .A1(reg_array_7__30_), .A2(n436), .B1(reg_array_6__30_), 
        .B2(n433), .C1(reg_array_5__30_), .C2(n430), .D1(reg_array_4__30_), 
        .D2(n427), .ZN(n478) );
  aoi2222d1 U474 ( .A1(reg_array_3__30_), .A2(n424), .B1(reg_array_2__30_), 
        .B2(n421), .C1(reg_array_1__30_), .C2(n418), .D1(reg_array_0__30_), 
        .D2(n404), .ZN(n479) );
  aoi2222d1 U475 ( .A1(test_so2), .A2(n436), .B1(reg_array_6__31_), .B2(n433), 
        .C1(reg_array_5__31_), .C2(n430), .D1(reg_array_4__31_), .D2(n427), 
        .ZN(n476) );
  aoi2222d1 U476 ( .A1(reg_array_3__31_), .A2(n424), .B1(reg_array_2__31_), 
        .B2(n421), .C1(reg_array_1__31_), .C2(n418), .D1(reg_array_0__31_), 
        .D2(n404), .ZN(n477) );
  nr03d0 U477 ( .A1(rd_addr_1_), .A2(rd_addr_2_), .A3(rd_addr_0_), .ZN(n538)
         );
  nr03d0 U478 ( .A1(rd_addr_1_), .A2(rd_addr_2_), .A3(n475), .ZN(n539) );
  nr03d0 U479 ( .A1(rd_addr_0_), .A2(rd_addr_2_), .A3(n474), .ZN(n540) );
  nr03d0 U480 ( .A1(n475), .A2(rd_addr_2_), .A3(n474), .ZN(n541) );
  nd04d0 U482 ( .A1(wr_addr_0_), .A2(n472), .A3(n471), .A4(n470), .ZN(n473) );
  nd04d0 U483 ( .A1(wr_addr_1_), .A2(n472), .A3(n468), .A4(n470), .ZN(n469) );
  nd04d0 U484 ( .A1(wr_addr_1_), .A2(wr_addr_0_), .A3(n472), .A4(n470), .ZN(
        n467) );
  nd04d0 U485 ( .A1(wr_addr_2_), .A2(n472), .A3(n468), .A4(n471), .ZN(n466) );
  nd04d0 U486 ( .A1(wr_addr_2_), .A2(wr_addr_0_), .A3(n472), .A4(n471), .ZN(
        n465) );
  nd04d0 U487 ( .A1(wr_addr_2_), .A2(wr_addr_1_), .A3(n472), .A4(n468), .ZN(
        n464) );
  nd04d0 U488 ( .A1(wr_addr_2_), .A2(wr_addr_1_), .A3(wr_addr_0_), .A4(n472), 
        .ZN(n463) );
  SDRAM_FIFO_1_DW_fifoctl_s2_sf_0 SD_FIFO_CTL ( .clk_push(fifo_clk_push), 
        .clk_pop(fifo_clk_pop), .rst_n(fifo_rst_n), .push_req_n(
        fifo_push_req_n), .pop_req_n(fifo_pop_req_n), .we_n(we_n), 
        .push_empty(push_empty_fifo), .push_ae(push_ae_fifo), .push_hf(
        push_hf_fifo), .push_af(push_af_fifo), .push_full(push_full_fifo), 
        .push_error(push_error_fifo), .pop_empty(pop_empty_fifo), .pop_ae(
        pop_ae_fifo), .pop_hf(pop_hf_fifo), .pop_af(pop_af_fifo), .pop_full(
        pop_full_fifo), .pop_error(pop_error_fifo), .wr_addr({wr_addr_2_, 
        wr_addr_1_, wr_addr_0_}), .rd_addr({rd_addr_2_, rd_addr_1_, rd_addr_0_}), .push_word_count({SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12}), .pop_word_count({
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16}), .test(test_mode), 
        .test_si1(test_si1), .test_si2(test_si2), .test_se(test_se), 
        .test_so2(n869), .test_so1(n872) );
  senrq1 reg_array_reg_0__31_ ( .D(N791), .SD(reg_array_0__30_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__31_) );
  senrq1 reg_array_reg_0__30_ ( .D(N789), .SD(reg_array_0__29_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__30_) );
  senrq1 reg_array_reg_0__29_ ( .D(N787), .SD(reg_array_0__28_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__29_) );
  senrq1 reg_array_reg_0__28_ ( .D(N785), .SD(reg_array_0__27_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__28_) );
  senrq1 reg_array_reg_0__27_ ( .D(N783), .SD(reg_array_0__26_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__27_) );
  senrq1 reg_array_reg_0__26_ ( .D(N781), .SD(reg_array_0__25_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__26_) );
  senrq1 reg_array_reg_0__25_ ( .D(N779), .SD(reg_array_0__24_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__25_) );
  senrq1 reg_array_reg_0__24_ ( .D(N777), .SD(reg_array_0__23_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__24_) );
  senrq1 reg_array_reg_0__23_ ( .D(N775), .SD(reg_array_0__22_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__23_) );
  senrq1 reg_array_reg_0__22_ ( .D(N773), .SD(reg_array_0__21_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__22_) );
  senrq1 reg_array_reg_0__21_ ( .D(N771), .SD(reg_array_0__20_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__21_) );
  senrq1 reg_array_reg_0__20_ ( .D(N769), .SD(reg_array_0__19_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__20_) );
  senrq1 reg_array_reg_0__19_ ( .D(N767), .SD(reg_array_0__18_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__19_) );
  senrq1 reg_array_reg_0__18_ ( .D(N765), .SD(reg_array_0__17_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__18_) );
  senrq1 reg_array_reg_0__17_ ( .D(N763), .SD(reg_array_0__16_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__17_) );
  senrq1 reg_array_reg_0__16_ ( .D(N761), .SD(reg_array_0__15_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__16_) );
  senrq1 reg_array_reg_0__15_ ( .D(N759), .SD(reg_array_0__14_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__15_) );
  senrq1 reg_array_reg_0__14_ ( .D(N757), .SD(reg_array_0__13_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__14_) );
  senrq1 reg_array_reg_0__13_ ( .D(N755), .SD(reg_array_0__12_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__13_) );
  senrq1 reg_array_reg_0__12_ ( .D(N753), .SD(reg_array_0__11_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__12_) );
  senrq1 reg_array_reg_0__11_ ( .D(N751), .SD(reg_array_0__10_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__11_) );
  senrq1 reg_array_reg_0__10_ ( .D(N749), .SD(reg_array_0__9_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__10_) );
  senrq1 reg_array_reg_0__9_ ( .D(N747), .SD(reg_array_0__8_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__9_) );
  senrq1 reg_array_reg_0__8_ ( .D(N745), .SD(reg_array_0__7_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__8_) );
  senrq1 reg_array_reg_0__7_ ( .D(N743), .SD(reg_array_0__6_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__7_) );
  senrq1 reg_array_reg_0__6_ ( .D(N741), .SD(reg_array_0__5_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__6_) );
  senrq1 reg_array_reg_0__5_ ( .D(N739), .SD(reg_array_0__4_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__5_) );
  senrq1 reg_array_reg_0__4_ ( .D(N737), .SD(reg_array_0__3_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__4_) );
  senrq1 reg_array_reg_0__3_ ( .D(N735), .SD(reg_array_0__2_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__3_) );
  senrq1 reg_array_reg_0__2_ ( .D(N733), .SD(reg_array_0__1_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__2_) );
  senrq1 reg_array_reg_0__1_ ( .D(N731), .SD(reg_array_0__0_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_0__1_) );
  senrq1 reg_array_reg_0__0_ ( .D(N729), .SD(n869), .ENN(n439), .SC(test_se), 
        .CP(fifo_clk_push), .Q(reg_array_0__0_) );
  senrq1 reg_array_reg_1__31_ ( .D(N791), .SD(reg_array_1__30_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__31_) );
  senrq1 reg_array_reg_1__30_ ( .D(N789), .SD(reg_array_1__29_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__30_) );
  senrq1 reg_array_reg_1__29_ ( .D(N787), .SD(reg_array_1__28_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__29_) );
  senrq1 reg_array_reg_1__28_ ( .D(N785), .SD(reg_array_1__27_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__28_) );
  senrq1 reg_array_reg_1__27_ ( .D(N783), .SD(reg_array_1__26_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__27_) );
  senrq1 reg_array_reg_1__26_ ( .D(N781), .SD(reg_array_1__25_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__26_) );
  senrq1 reg_array_reg_1__25_ ( .D(N779), .SD(reg_array_1__24_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__25_) );
  senrq1 reg_array_reg_1__24_ ( .D(N777), .SD(reg_array_1__23_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__24_) );
  senrq1 reg_array_reg_1__23_ ( .D(N775), .SD(reg_array_1__22_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__23_) );
  senrq1 reg_array_reg_1__22_ ( .D(N773), .SD(reg_array_1__21_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__22_) );
  senrq1 reg_array_reg_1__21_ ( .D(N771), .SD(reg_array_1__20_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__21_) );
  senrq1 reg_array_reg_1__20_ ( .D(N769), .SD(reg_array_1__19_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__20_) );
  senrq1 reg_array_reg_1__19_ ( .D(N767), .SD(reg_array_1__18_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__19_) );
  senrq1 reg_array_reg_1__18_ ( .D(N765), .SD(reg_array_1__17_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__18_) );
  senrq1 reg_array_reg_1__17_ ( .D(N763), .SD(reg_array_1__16_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__17_) );
  senrq1 reg_array_reg_1__16_ ( .D(N761), .SD(reg_array_1__15_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__16_) );
  senrq1 reg_array_reg_1__15_ ( .D(N759), .SD(reg_array_1__14_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__15_) );
  senrq1 reg_array_reg_1__14_ ( .D(N757), .SD(reg_array_1__13_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__14_) );
  senrq1 reg_array_reg_1__13_ ( .D(N755), .SD(reg_array_1__12_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__13_) );
  senrq1 reg_array_reg_1__12_ ( .D(N753), .SD(reg_array_1__11_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__12_) );
  senrq1 reg_array_reg_1__11_ ( .D(N751), .SD(reg_array_1__10_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__11_) );
  senrq1 reg_array_reg_1__10_ ( .D(N749), .SD(reg_array_1__9_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__10_) );
  senrq1 reg_array_reg_1__9_ ( .D(N747), .SD(reg_array_1__8_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__9_) );
  senrq1 reg_array_reg_1__8_ ( .D(N745), .SD(reg_array_1__7_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__8_) );
  senrq1 reg_array_reg_1__7_ ( .D(N743), .SD(reg_array_1__6_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__7_) );
  senrq1 reg_array_reg_1__6_ ( .D(N741), .SD(reg_array_1__5_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__6_) );
  senrq1 reg_array_reg_1__5_ ( .D(N739), .SD(reg_array_1__4_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__5_) );
  senrq1 reg_array_reg_1__4_ ( .D(N737), .SD(reg_array_1__3_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__4_) );
  senrq1 reg_array_reg_1__3_ ( .D(N735), .SD(reg_array_1__2_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__3_) );
  senrq1 reg_array_reg_1__2_ ( .D(N733), .SD(reg_array_1__1_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__2_) );
  senrq1 reg_array_reg_1__1_ ( .D(N731), .SD(reg_array_1__0_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__1_) );
  senrq1 reg_array_reg_1__0_ ( .D(N729), .SD(reg_array_0__31_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_1__0_) );
  senrq1 reg_array_reg_2__31_ ( .D(N791), .SD(reg_array_2__30_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__31_) );
  senrq1 reg_array_reg_2__30_ ( .D(N789), .SD(reg_array_2__29_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__30_) );
  senrq1 reg_array_reg_2__29_ ( .D(N787), .SD(reg_array_2__28_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__29_) );
  senrq1 reg_array_reg_2__28_ ( .D(N785), .SD(reg_array_2__27_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__28_) );
  senrq1 reg_array_reg_2__27_ ( .D(N783), .SD(reg_array_2__26_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__27_) );
  senrq1 reg_array_reg_2__26_ ( .D(N781), .SD(reg_array_2__25_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__26_) );
  senrq1 reg_array_reg_2__25_ ( .D(N779), .SD(reg_array_2__24_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__25_) );
  senrq1 reg_array_reg_2__24_ ( .D(N777), .SD(reg_array_2__23_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__24_) );
  senrq1 reg_array_reg_2__23_ ( .D(N775), .SD(reg_array_2__22_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__23_) );
  senrq1 reg_array_reg_2__22_ ( .D(N773), .SD(reg_array_2__21_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__22_) );
  senrq1 reg_array_reg_2__21_ ( .D(N771), .SD(reg_array_2__20_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__21_) );
  senrq1 reg_array_reg_2__20_ ( .D(N769), .SD(reg_array_2__19_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__20_) );
  senrq1 reg_array_reg_2__19_ ( .D(N767), .SD(reg_array_2__18_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__19_) );
  senrq1 reg_array_reg_2__18_ ( .D(N765), .SD(reg_array_2__17_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__18_) );
  senrq1 reg_array_reg_2__17_ ( .D(N763), .SD(reg_array_2__16_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__17_) );
  senrq1 reg_array_reg_2__16_ ( .D(N761), .SD(reg_array_2__15_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__16_) );
  senrq1 reg_array_reg_2__15_ ( .D(N759), .SD(reg_array_2__14_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__15_) );
  senrq1 reg_array_reg_2__14_ ( .D(N757), .SD(reg_array_2__13_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__14_) );
  senrq1 reg_array_reg_2__13_ ( .D(N755), .SD(reg_array_2__12_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__13_) );
  senrq1 reg_array_reg_2__12_ ( .D(N753), .SD(reg_array_2__11_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__12_) );
  senrq1 reg_array_reg_2__11_ ( .D(N751), .SD(reg_array_2__10_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__11_) );
  senrq1 reg_array_reg_2__10_ ( .D(N749), .SD(reg_array_2__9_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__10_) );
  senrq1 reg_array_reg_2__9_ ( .D(N747), .SD(reg_array_2__8_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__9_) );
  senrq1 reg_array_reg_2__8_ ( .D(N745), .SD(reg_array_2__7_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__8_) );
  senrq1 reg_array_reg_2__7_ ( .D(N743), .SD(reg_array_2__6_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__7_) );
  senrq1 reg_array_reg_2__6_ ( .D(N741), .SD(reg_array_2__5_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__6_) );
  senrq1 reg_array_reg_2__5_ ( .D(N739), .SD(reg_array_2__4_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__5_) );
  senrq1 reg_array_reg_2__4_ ( .D(N737), .SD(reg_array_2__3_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__4_) );
  senrq1 reg_array_reg_2__3_ ( .D(N735), .SD(reg_array_2__2_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__3_) );
  senrq1 reg_array_reg_2__2_ ( .D(N733), .SD(reg_array_2__1_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__2_) );
  senrq1 reg_array_reg_2__1_ ( .D(N731), .SD(reg_array_2__0_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__1_) );
  senrq1 reg_array_reg_2__0_ ( .D(N729), .SD(reg_array_1__31_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_2__0_) );
  senrq1 reg_array_reg_3__31_ ( .D(N791), .SD(reg_array_3__30_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__31_) );
  senrq1 reg_array_reg_3__30_ ( .D(N789), .SD(reg_array_3__29_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__30_) );
  senrq1 reg_array_reg_3__29_ ( .D(N787), .SD(reg_array_3__28_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__29_) );
  senrq1 reg_array_reg_3__28_ ( .D(N785), .SD(reg_array_3__27_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__28_) );
  senrq1 reg_array_reg_3__27_ ( .D(N783), .SD(reg_array_3__26_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__27_) );
  senrq1 reg_array_reg_3__26_ ( .D(N781), .SD(reg_array_3__25_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__26_) );
  senrq1 reg_array_reg_3__25_ ( .D(N779), .SD(reg_array_3__24_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__25_) );
  senrq1 reg_array_reg_3__24_ ( .D(N777), .SD(reg_array_3__23_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__24_) );
  senrq1 reg_array_reg_3__23_ ( .D(N775), .SD(reg_array_3__22_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__23_) );
  senrq1 reg_array_reg_3__22_ ( .D(N773), .SD(reg_array_3__21_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__22_) );
  senrq1 reg_array_reg_3__21_ ( .D(N771), .SD(reg_array_3__20_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__21_) );
  senrq1 reg_array_reg_3__20_ ( .D(N769), .SD(reg_array_3__19_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__20_) );
  senrq1 reg_array_reg_3__19_ ( .D(N767), .SD(reg_array_3__18_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__19_) );
  senrq1 reg_array_reg_3__18_ ( .D(N765), .SD(reg_array_3__17_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__18_) );
  senrq1 reg_array_reg_3__17_ ( .D(N763), .SD(reg_array_3__16_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__17_) );
  senrq1 reg_array_reg_3__16_ ( .D(N761), .SD(reg_array_3__15_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__16_) );
  senrq1 reg_array_reg_3__15_ ( .D(N759), .SD(reg_array_3__14_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__15_) );
  senrq1 reg_array_reg_3__14_ ( .D(N757), .SD(reg_array_3__13_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__14_) );
  senrq1 reg_array_reg_3__13_ ( .D(N755), .SD(reg_array_3__12_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__13_) );
  senrq1 reg_array_reg_3__12_ ( .D(N753), .SD(reg_array_3__11_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__12_) );
  senrq1 reg_array_reg_3__11_ ( .D(N751), .SD(reg_array_3__10_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__11_) );
  senrq1 reg_array_reg_3__10_ ( .D(N749), .SD(reg_array_3__9_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__10_) );
  senrq1 reg_array_reg_3__9_ ( .D(N747), .SD(reg_array_3__8_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__9_) );
  senrq1 reg_array_reg_3__8_ ( .D(N745), .SD(reg_array_3__7_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__8_) );
  senrq1 reg_array_reg_3__7_ ( .D(N743), .SD(reg_array_3__6_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__7_) );
  senrq1 reg_array_reg_3__6_ ( .D(N741), .SD(reg_array_3__5_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__6_) );
  senrq1 reg_array_reg_3__5_ ( .D(N739), .SD(reg_array_3__4_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__5_) );
  senrq1 reg_array_reg_3__4_ ( .D(N737), .SD(reg_array_3__3_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__4_) );
  senrq1 reg_array_reg_3__3_ ( .D(N735), .SD(reg_array_3__2_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__3_) );
  senrq1 reg_array_reg_3__2_ ( .D(N733), .SD(reg_array_3__1_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__2_) );
  senrq1 reg_array_reg_3__1_ ( .D(N731), .SD(reg_array_3__0_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__1_) );
  senrq1 reg_array_reg_3__0_ ( .D(N729), .SD(reg_array_2__31_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_3__0_) );
  senrq1 reg_array_reg_4__31_ ( .D(N791), .SD(reg_array_4__30_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__31_) );
  senrq1 reg_array_reg_4__30_ ( .D(N789), .SD(reg_array_4__29_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__30_) );
  senrq1 reg_array_reg_4__29_ ( .D(N787), .SD(reg_array_4__28_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__29_) );
  senrq1 reg_array_reg_4__28_ ( .D(N785), .SD(reg_array_4__27_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__28_) );
  senrq1 reg_array_reg_4__27_ ( .D(N783), .SD(reg_array_4__26_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__27_) );
  senrq1 reg_array_reg_4__26_ ( .D(N781), .SD(reg_array_4__25_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__26_) );
  senrq1 reg_array_reg_4__25_ ( .D(N779), .SD(reg_array_4__24_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__25_) );
  senrq1 reg_array_reg_4__24_ ( .D(N777), .SD(reg_array_4__23_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__24_) );
  senrq1 reg_array_reg_4__23_ ( .D(N775), .SD(reg_array_4__22_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__23_) );
  senrq1 reg_array_reg_4__22_ ( .D(N773), .SD(reg_array_4__21_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__22_) );
  senrq1 reg_array_reg_4__21_ ( .D(N771), .SD(reg_array_4__20_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__21_) );
  senrq1 reg_array_reg_4__20_ ( .D(N769), .SD(reg_array_4__19_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__20_) );
  senrq1 reg_array_reg_4__19_ ( .D(N767), .SD(reg_array_4__18_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__19_) );
  senrq1 reg_array_reg_4__18_ ( .D(N765), .SD(reg_array_4__17_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__18_) );
  senrq1 reg_array_reg_4__17_ ( .D(N763), .SD(reg_array_4__16_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__17_) );
  senrq1 reg_array_reg_4__16_ ( .D(N761), .SD(reg_array_4__15_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__16_) );
  senrq1 reg_array_reg_4__15_ ( .D(N759), .SD(reg_array_4__14_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__15_) );
  senrq1 reg_array_reg_4__14_ ( .D(N757), .SD(reg_array_4__13_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__14_) );
  senrq1 reg_array_reg_4__13_ ( .D(N755), .SD(reg_array_4__12_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__13_) );
  senrq1 reg_array_reg_4__12_ ( .D(N753), .SD(reg_array_4__11_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__12_) );
  senrq1 reg_array_reg_4__11_ ( .D(N751), .SD(reg_array_4__10_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__11_) );
  senrq1 reg_array_reg_4__10_ ( .D(N749), .SD(reg_array_4__9_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__10_) );
  senrq1 reg_array_reg_4__9_ ( .D(N747), .SD(reg_array_4__8_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__9_) );
  senrq1 reg_array_reg_4__8_ ( .D(N745), .SD(reg_array_4__7_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__8_) );
  senrq1 reg_array_reg_4__7_ ( .D(N743), .SD(reg_array_4__6_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__7_) );
  senrq1 reg_array_reg_4__6_ ( .D(N741), .SD(reg_array_4__5_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__6_) );
  senrq1 reg_array_reg_4__5_ ( .D(N739), .SD(reg_array_4__4_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__5_) );
  senrq1 reg_array_reg_4__4_ ( .D(N737), .SD(reg_array_4__3_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__4_) );
  senrq1 reg_array_reg_4__3_ ( .D(N735), .SD(reg_array_4__2_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__3_) );
  senrq1 reg_array_reg_4__2_ ( .D(N733), .SD(reg_array_4__1_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__2_) );
  senrq1 reg_array_reg_4__1_ ( .D(N731), .SD(reg_array_4__0_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__1_) );
  senrq1 reg_array_reg_4__0_ ( .D(N729), .SD(reg_array_3__31_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_4__0_) );
  senrq1 reg_array_reg_5__31_ ( .D(N791), .SD(reg_array_5__30_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__31_) );
  senrq1 reg_array_reg_5__30_ ( .D(N789), .SD(reg_array_5__29_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__30_) );
  senrq1 reg_array_reg_5__29_ ( .D(N787), .SD(reg_array_5__28_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__29_) );
  senrq1 reg_array_reg_5__28_ ( .D(N785), .SD(reg_array_5__27_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__28_) );
  senrq1 reg_array_reg_5__27_ ( .D(N783), .SD(reg_array_5__26_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__27_) );
  senrq1 reg_array_reg_5__26_ ( .D(N781), .SD(reg_array_5__25_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__26_) );
  senrq1 reg_array_reg_5__25_ ( .D(N779), .SD(reg_array_5__24_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__25_) );
  senrq1 reg_array_reg_5__24_ ( .D(N777), .SD(reg_array_5__23_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__24_) );
  senrq1 reg_array_reg_5__23_ ( .D(N775), .SD(reg_array_5__22_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__23_) );
  senrq1 reg_array_reg_5__22_ ( .D(N773), .SD(reg_array_5__21_), .ENN(n456), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__22_) );
  senrq1 reg_array_reg_5__21_ ( .D(N771), .SD(reg_array_5__20_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__21_) );
  senrq1 reg_array_reg_5__20_ ( .D(N769), .SD(reg_array_5__19_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__20_) );
  senrq1 reg_array_reg_5__19_ ( .D(N767), .SD(reg_array_5__18_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__19_) );
  senrq1 reg_array_reg_5__18_ ( .D(N765), .SD(reg_array_5__17_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__18_) );
  senrq1 reg_array_reg_5__17_ ( .D(N763), .SD(reg_array_5__16_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__17_) );
  senrq1 reg_array_reg_5__16_ ( .D(N761), .SD(reg_array_5__15_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__16_) );
  senrq1 reg_array_reg_5__15_ ( .D(N759), .SD(reg_array_5__14_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__15_) );
  senrq1 reg_array_reg_5__14_ ( .D(N757), .SD(reg_array_5__13_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__14_) );
  senrq1 reg_array_reg_5__13_ ( .D(N755), .SD(reg_array_5__12_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__13_) );
  senrq1 reg_array_reg_5__12_ ( .D(N753), .SD(reg_array_5__11_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__12_) );
  senrq1 reg_array_reg_5__11_ ( .D(N751), .SD(reg_array_5__10_), .ENN(n455), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__11_) );
  senrq1 reg_array_reg_5__10_ ( .D(N749), .SD(reg_array_5__9_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__10_) );
  senrq1 reg_array_reg_5__9_ ( .D(N747), .SD(reg_array_5__8_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__9_) );
  senrq1 reg_array_reg_5__8_ ( .D(N745), .SD(reg_array_5__7_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__8_) );
  senrq1 reg_array_reg_5__7_ ( .D(N743), .SD(reg_array_5__6_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__7_) );
  senrq1 reg_array_reg_5__6_ ( .D(N741), .SD(reg_array_5__5_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__6_) );
  senrq1 reg_array_reg_5__5_ ( .D(N739), .SD(reg_array_5__4_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__5_) );
  senrq1 reg_array_reg_5__4_ ( .D(N737), .SD(reg_array_5__3_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__4_) );
  senrq1 reg_array_reg_5__3_ ( .D(N735), .SD(reg_array_5__2_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__3_) );
  senrq1 reg_array_reg_5__2_ ( .D(N733), .SD(reg_array_5__1_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__2_) );
  senrq1 reg_array_reg_5__1_ ( .D(N731), .SD(reg_array_5__0_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__1_) );
  senrq1 reg_array_reg_5__0_ ( .D(N729), .SD(reg_array_4__31_), .ENN(n454), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_5__0_) );
  senrq1 reg_array_reg_6__31_ ( .D(N791), .SD(reg_array_6__30_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__31_) );
  senrq1 reg_array_reg_6__30_ ( .D(N789), .SD(reg_array_6__29_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__30_) );
  senrq1 reg_array_reg_6__29_ ( .D(N787), .SD(reg_array_6__28_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__29_) );
  senrq1 reg_array_reg_6__28_ ( .D(N785), .SD(reg_array_6__27_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__28_) );
  senrq1 reg_array_reg_6__27_ ( .D(N783), .SD(reg_array_6__26_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__27_) );
  senrq1 reg_array_reg_6__26_ ( .D(N781), .SD(reg_array_6__25_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__26_) );
  senrq1 reg_array_reg_6__25_ ( .D(N779), .SD(reg_array_6__24_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__25_) );
  senrq1 reg_array_reg_6__24_ ( .D(N777), .SD(reg_array_6__23_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__24_) );
  senrq1 reg_array_reg_6__23_ ( .D(N775), .SD(reg_array_6__22_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__23_) );
  senrq1 reg_array_reg_6__22_ ( .D(N773), .SD(reg_array_6__21_), .ENN(n459), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__22_) );
  senrq1 reg_array_reg_6__21_ ( .D(N771), .SD(reg_array_6__20_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__21_) );
  senrq1 reg_array_reg_6__20_ ( .D(N769), .SD(reg_array_6__19_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__20_) );
  senrq1 reg_array_reg_6__19_ ( .D(N767), .SD(reg_array_6__18_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__19_) );
  senrq1 reg_array_reg_6__18_ ( .D(N765), .SD(reg_array_6__17_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__18_) );
  senrq1 reg_array_reg_6__17_ ( .D(N763), .SD(reg_array_6__16_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__17_) );
  senrq1 reg_array_reg_6__16_ ( .D(N761), .SD(reg_array_6__15_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__16_) );
  senrq1 reg_array_reg_6__15_ ( .D(N759), .SD(reg_array_6__14_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__15_) );
  senrq1 reg_array_reg_6__14_ ( .D(N757), .SD(reg_array_6__13_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__14_) );
  senrq1 reg_array_reg_6__13_ ( .D(N755), .SD(reg_array_6__12_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__13_) );
  senrq1 reg_array_reg_6__12_ ( .D(N753), .SD(reg_array_6__11_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__12_) );
  senrq1 reg_array_reg_6__11_ ( .D(N751), .SD(reg_array_6__10_), .ENN(n458), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__11_) );
  senrq1 reg_array_reg_6__10_ ( .D(N749), .SD(reg_array_6__9_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__10_) );
  senrq1 reg_array_reg_6__9_ ( .D(N747), .SD(reg_array_6__8_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__9_) );
  senrq1 reg_array_reg_6__8_ ( .D(N745), .SD(reg_array_6__7_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__8_) );
  senrq1 reg_array_reg_6__7_ ( .D(N743), .SD(reg_array_6__6_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__7_) );
  senrq1 reg_array_reg_6__6_ ( .D(N741), .SD(reg_array_6__5_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__6_) );
  senrq1 reg_array_reg_6__5_ ( .D(N739), .SD(reg_array_6__4_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__5_) );
  senrq1 reg_array_reg_6__4_ ( .D(N737), .SD(reg_array_6__3_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__4_) );
  senrq1 reg_array_reg_6__3_ ( .D(N735), .SD(reg_array_6__2_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__3_) );
  senrq1 reg_array_reg_6__2_ ( .D(N733), .SD(reg_array_6__1_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__2_) );
  senrq1 reg_array_reg_6__1_ ( .D(N731), .SD(reg_array_6__0_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__1_) );
  senrq1 reg_array_reg_6__0_ ( .D(N729), .SD(reg_array_5__31_), .ENN(n457), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_6__0_) );
  senrq1 reg_array_reg_7__31_ ( .D(N791), .SD(reg_array_7__30_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(test_so2) );
  senrq1 reg_array_reg_7__30_ ( .D(N789), .SD(reg_array_7__29_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__30_) );
  senrq1 reg_array_reg_7__29_ ( .D(N787), .SD(reg_array_7__28_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__29_) );
  senrq1 reg_array_reg_7__28_ ( .D(N785), .SD(reg_array_7__27_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__28_) );
  senrq1 reg_array_reg_7__27_ ( .D(N783), .SD(reg_array_7__26_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__27_) );
  senrq1 reg_array_reg_7__26_ ( .D(N781), .SD(reg_array_7__25_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__26_) );
  senrq1 reg_array_reg_7__25_ ( .D(N779), .SD(reg_array_7__24_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__25_) );
  senrq1 reg_array_reg_7__24_ ( .D(N777), .SD(reg_array_7__23_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__24_) );
  senrq1 reg_array_reg_7__23_ ( .D(N775), .SD(reg_array_7__22_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__23_) );
  senrq1 reg_array_reg_7__22_ ( .D(N773), .SD(reg_array_7__21_), .ENN(n462), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__22_) );
  senrq1 reg_array_reg_7__21_ ( .D(N771), .SD(reg_array_7__20_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__21_) );
  senrq1 reg_array_reg_7__20_ ( .D(N769), .SD(reg_array_7__19_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__20_) );
  senrq1 reg_array_reg_7__19_ ( .D(N767), .SD(reg_array_7__18_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__19_) );
  senrq1 reg_array_reg_7__18_ ( .D(N765), .SD(reg_array_7__17_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__18_) );
  senrq1 reg_array_reg_7__17_ ( .D(N763), .SD(reg_array_7__16_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__17_) );
  senrq1 reg_array_reg_7__16_ ( .D(N761), .SD(reg_array_7__15_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__16_) );
  senrq1 reg_array_reg_7__15_ ( .D(N759), .SD(reg_array_7__14_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__15_) );
  senrq1 reg_array_reg_7__14_ ( .D(N757), .SD(reg_array_7__13_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__14_) );
  senrq1 reg_array_reg_7__13_ ( .D(N755), .SD(reg_array_7__12_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__13_) );
  senrq1 reg_array_reg_7__12_ ( .D(N753), .SD(reg_array_7__11_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__12_) );
  senrq1 reg_array_reg_7__11_ ( .D(N751), .SD(reg_array_7__10_), .ENN(n461), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__11_) );
  senrq1 reg_array_reg_7__10_ ( .D(N749), .SD(reg_array_7__9_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__10_) );
  senrq1 reg_array_reg_7__9_ ( .D(N747), .SD(reg_array_7__8_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__9_) );
  senrq1 reg_array_reg_7__8_ ( .D(N745), .SD(reg_array_7__7_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__8_) );
  senrq1 reg_array_reg_7__7_ ( .D(N743), .SD(reg_array_7__6_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__7_) );
  senrq1 reg_array_reg_7__6_ ( .D(N741), .SD(reg_array_7__5_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__6_) );
  senrq1 reg_array_reg_7__5_ ( .D(N739), .SD(reg_array_7__4_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__5_) );
  senrq1 reg_array_reg_7__4_ ( .D(N737), .SD(reg_array_7__3_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__4_) );
  senrq1 reg_array_reg_7__3_ ( .D(N735), .SD(reg_array_7__2_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__3_) );
  senrq1 reg_array_reg_7__2_ ( .D(N733), .SD(reg_array_7__1_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__2_) );
  senrq1 reg_array_reg_7__1_ ( .D(N731), .SD(reg_array_7__0_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__1_) );
  senrq1 reg_array_reg_7__0_ ( .D(N729), .SD(reg_array_6__31_), .ENN(n460), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_7__0_) );
  sdnrq1 data_out_sync_reg_31_ ( .D(N807), .SD(data_out_sync_30_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_31_) );
  sdnrq1 data_out_sync_reg_30_ ( .D(N808), .SD(data_out_sync_29_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_30_) );
  sdnrq1 data_out_sync_reg_29_ ( .D(N809), .SD(data_out_sync_28_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_29_) );
  sdnrq1 data_out_sync_reg_28_ ( .D(N810), .SD(data_out_sync_27_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_28_) );
  sdnrq1 data_out_sync_reg_27_ ( .D(N811), .SD(data_out_sync_26_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_27_) );
  sdnrq1 data_out_sync_reg_26_ ( .D(N812), .SD(data_out_sync_25_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_26_) );
  sdnrq1 data_out_sync_reg_25_ ( .D(N813), .SD(data_out_sync_24_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_25_) );
  sdnrq1 data_out_sync_reg_24_ ( .D(N814), .SD(data_out_sync_23_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_24_) );
  sdnrq1 data_out_sync_reg_23_ ( .D(N815), .SD(data_out_sync_22_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_23_) );
  sdnrq1 data_out_sync_reg_22_ ( .D(N816), .SD(data_out_sync_21_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_22_) );
  sdnrq1 data_out_sync_reg_21_ ( .D(N817), .SD(data_out_sync_20_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_21_) );
  sdnrq1 data_out_sync_reg_20_ ( .D(N818), .SD(data_out_sync_19_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_20_) );
  sdnrq1 data_out_sync_reg_19_ ( .D(N819), .SD(data_out_sync_18_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_19_) );
  sdnrq1 data_out_sync_reg_18_ ( .D(N820), .SD(data_out_sync_17_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_18_) );
  sdnrq1 data_out_sync_reg_17_ ( .D(N821), .SD(data_out_sync_16_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_17_) );
  sdnrq1 data_out_sync_reg_16_ ( .D(N822), .SD(data_out_sync_15_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_16_) );
  sdnrq1 data_out_sync_reg_15_ ( .D(N823), .SD(data_out_sync_14_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_15_) );
  sdnrq1 data_out_sync_reg_14_ ( .D(N824), .SD(data_out_sync_13_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_14_) );
  sdnrq1 data_out_sync_reg_13_ ( .D(N825), .SD(data_out_sync_12_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_13_) );
  sdnrq1 data_out_sync_reg_12_ ( .D(N826), .SD(data_out_sync_11_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_12_) );
  sdnrq1 data_out_sync_reg_11_ ( .D(N827), .SD(data_out_sync_10_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_11_) );
  sdnrq1 data_out_sync_reg_10_ ( .D(N828), .SD(data_out_sync_9_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_10_) );
  sdnrq1 data_out_sync_reg_9_ ( .D(N829), .SD(data_out_sync_8_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_9_) );
  sdnrq1 data_out_sync_reg_8_ ( .D(N830), .SD(data_out_sync_7_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_8_) );
  sdnrq1 data_out_sync_reg_7_ ( .D(N831), .SD(data_out_sync_6_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_7_) );
  sdnrq1 data_out_sync_reg_6_ ( .D(N832), .SD(data_out_sync_5_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_6_) );
  sdnrq1 data_out_sync_reg_5_ ( .D(N833), .SD(data_out_sync_4_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_5_) );
  sdnrq1 data_out_sync_reg_4_ ( .D(N834), .SD(data_out_sync_3_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_4_) );
  sdnrq1 data_out_sync_reg_3_ ( .D(N835), .SD(data_out_sync_2_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_3_) );
  sdnrq1 data_out_sync_reg_2_ ( .D(N836), .SD(data_out_sync_1_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_2_) );
  sdnrq1 data_out_sync_reg_1_ ( .D(N837), .SD(data_out_sync_0_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_1_) );
  sdnrq1 data_out_sync_reg_0_ ( .D(N838), .SD(data_out_fifo[31]), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_0_) );
  sdnrq1 data_out_reg_15_ ( .D(data_out_sync_15_), .SD(data_out_fifo[14]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[15]) );
  sdnrq1 data_out_reg_14_ ( .D(data_out_sync_14_), .SD(data_out_fifo[13]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[14]) );
  sdnrq1 data_out_reg_13_ ( .D(data_out_sync_13_), .SD(data_out_fifo[12]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[13]) );
  sdnrq1 data_out_reg_12_ ( .D(data_out_sync_12_), .SD(data_out_fifo[11]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[12]) );
  sdnrq1 data_out_reg_11_ ( .D(data_out_sync_11_), .SD(data_out_fifo[10]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[11]) );
  sdnrq1 data_out_reg_10_ ( .D(data_out_sync_10_), .SD(data_out_fifo[9]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[10]) );
  sdnrq1 data_out_reg_9_ ( .D(data_out_sync_9_), .SD(data_out_fifo[8]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[9]) );
  sdnrq1 data_out_reg_8_ ( .D(data_out_sync_8_), .SD(data_out_fifo[7]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[8]) );
  sdnrq1 data_out_reg_7_ ( .D(data_out_sync_7_), .SD(data_out_fifo[6]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[7]) );
  sdnrq1 data_out_reg_6_ ( .D(data_out_sync_6_), .SD(data_out_fifo[5]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[6]) );
  sdnrq1 data_out_reg_5_ ( .D(data_out_sync_5_), .SD(data_out_fifo[4]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[5]) );
  sdnrq1 data_out_reg_4_ ( .D(data_out_sync_4_), .SD(data_out_fifo[3]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[4]) );
  sdnrq1 data_out_reg_3_ ( .D(data_out_sync_3_), .SD(data_out_fifo[2]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[3]) );
  sdnrq1 data_out_reg_2_ ( .D(data_out_sync_2_), .SD(data_out_fifo[1]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[2]) );
  sdnrq1 data_out_reg_1_ ( .D(data_out_sync_1_), .SD(data_out_fifo[0]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[1]) );
  sdnrq1 data_out_reg_0_ ( .D(data_out_sync_0_), .SD(n872), .SC(test_se), .CP(
        fifo_clk_pop), .Q(data_out_fifo[0]) );
  sdnrq1 data_out_reg_31_ ( .D(data_out_sync_31_), .SD(data_out_fifo[30]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[31]) );
  sdnrq1 data_out_reg_30_ ( .D(data_out_sync_30_), .SD(data_out_fifo[29]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[30]) );
  sdnrq1 data_out_reg_29_ ( .D(data_out_sync_29_), .SD(data_out_fifo[28]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[29]) );
  sdnrq1 data_out_reg_28_ ( .D(data_out_sync_28_), .SD(data_out_fifo[27]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[28]) );
  sdnrq1 data_out_reg_27_ ( .D(data_out_sync_27_), .SD(data_out_fifo[26]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[27]) );
  sdnrq1 data_out_reg_26_ ( .D(data_out_sync_26_), .SD(data_out_fifo[25]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[26]) );
  sdnrq1 data_out_reg_25_ ( .D(data_out_sync_25_), .SD(data_out_fifo[24]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[25]) );
  sdnrq1 data_out_reg_24_ ( .D(data_out_sync_24_), .SD(data_out_fifo[23]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[24]) );
  sdnrq1 data_out_reg_23_ ( .D(data_out_sync_23_), .SD(data_out_fifo[22]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[23]) );
  sdnrq1 data_out_reg_22_ ( .D(data_out_sync_22_), .SD(data_out_fifo[21]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[22]) );
  sdnrq1 data_out_reg_21_ ( .D(data_out_sync_21_), .SD(data_out_fifo[20]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[21]) );
  sdnrq1 data_out_reg_20_ ( .D(data_out_sync_20_), .SD(data_out_fifo[19]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[20]) );
  sdnrq1 data_out_reg_19_ ( .D(data_out_sync_19_), .SD(data_out_fifo[18]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[19]) );
  sdnrq1 data_out_reg_18_ ( .D(data_out_sync_18_), .SD(data_out_fifo[17]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[18]) );
  sdnrq1 data_out_reg_17_ ( .D(data_out_sync_17_), .SD(data_out_fifo[16]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[17]) );
  sdnrq1 data_out_reg_16_ ( .D(data_out_sync_16_), .SD(data_out_fifo[15]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[16]) );
  inv0d1 U98 ( .I(we_n), .ZN(n472) );
  bufbd1 U131 ( .I(n540), .Z(n422) );
  bufbd1 U164 ( .I(n538), .Z(n416) );
  bufbd1 U197 ( .I(n541), .Z(n425) );
  bufbd1 U230 ( .I(n539), .Z(n419) );
  bufbd1 U263 ( .I(n540), .Z(n421) );
  bufbd1 U296 ( .I(n538), .Z(n404) );
  bufbd1 U329 ( .I(n541), .Z(n424) );
  bufbd1 U331 ( .I(n539), .Z(n418) );
  bufbd1 U332 ( .I(n130), .Z(n460) );
  bufbd1 U333 ( .I(n130), .Z(n461) );
  bufbd1 U334 ( .I(n1), .Z(n457) );
  bufbd1 U335 ( .I(n1), .Z(n458) );
  bufbd1 U336 ( .I(n97), .Z(n454) );
  bufbd1 U337 ( .I(n97), .Z(n455) );
  bufbd1 U338 ( .I(n229), .Z(n451) );
  bufbd1 U339 ( .I(n229), .Z(n452) );
  bufbd1 U340 ( .I(n163), .Z(n448) );
  bufbd1 U341 ( .I(n163), .Z(n449) );
  bufbd1 U342 ( .I(n196), .Z(n445) );
  bufbd1 U343 ( .I(n196), .Z(n446) );
  bufbd1 U344 ( .I(n262), .Z(n442) );
  bufbd1 U345 ( .I(n262), .Z(n443) );
  bufbd1 U346 ( .I(n295), .Z(n439) );
  bufbd1 U347 ( .I(n295), .Z(n440) );
  bufbd1 U348 ( .I(n540), .Z(n423) );
  bufbd1 U349 ( .I(n538), .Z(n417) );
  bufbd1 U350 ( .I(n541), .Z(n426) );
  bufbd1 U351 ( .I(n539), .Z(n420) );
  bufbd1 U352 ( .I(n130), .Z(n462) );
  bufbd1 U353 ( .I(n1), .Z(n459) );
  bufbd1 U354 ( .I(n97), .Z(n456) );
  bufbd1 U355 ( .I(n229), .Z(n453) );
  bufbd1 U356 ( .I(n163), .Z(n450) );
  bufbd1 U357 ( .I(n196), .Z(n447) );
  bufbd1 U358 ( .I(n262), .Z(n444) );
  bufbd1 U359 ( .I(n295), .Z(n441) );
  bufbd1 U360 ( .I(n544), .Z(n434) );
  bufbd1 U361 ( .I(n542), .Z(n428) );
  bufbd1 U362 ( .I(n543), .Z(n431) );
  bufbd1 U367 ( .I(n545), .Z(n437) );
  bufbd1 U368 ( .I(n544), .Z(n433) );
  bufbd1 U369 ( .I(n542), .Z(n427) );
  bufbd1 U370 ( .I(n543), .Z(n430) );
  bufbd1 U371 ( .I(n545), .Z(n436) );
  bufbd1 U372 ( .I(n544), .Z(n435) );
  bufbd1 U373 ( .I(n542), .Z(n429) );
  bufbd1 U374 ( .I(n543), .Z(n432) );
  bufbd1 U375 ( .I(n545), .Z(n438) );
  an02d1 U376 ( .A1(fifo_rst_n), .A2(n464), .Z(n1) );
  an02d1 U377 ( .A1(fifo_rst_n), .A2(n465), .Z(n97) );
  inv0d1 U378 ( .I(rd_addr_1_), .ZN(n474) );
  inv0d1 U411 ( .I(rd_addr_0_), .ZN(n475) );
  an02d1 U412 ( .A1(fifo_rst_n), .A2(n463), .Z(n130) );
  an02d1 U481 ( .A1(fifo_rst_n), .A2(n467), .Z(n163) );
  an02d1 U489 ( .A1(fifo_rst_n), .A2(n469), .Z(n196) );
  an02d1 U490 ( .A1(fifo_rst_n), .A2(n466), .Z(n229) );
  an02d1 U491 ( .A1(fifo_rst_n), .A2(n473), .Z(n262) );
  an02d1 U492 ( .A1(n328), .A2(fifo_rst_n), .Z(n295) );
  or04d1 U493 ( .A1(wr_addr_2_), .A2(wr_addr_1_), .A3(wr_addr_0_), .A4(we_n), 
        .Z(n328) );
  nd02d1 U494 ( .A1(n547), .A2(n546), .ZN(N838) );
  nd02d1 U495 ( .A1(n537), .A2(n536), .ZN(N837) );
  nd02d1 U496 ( .A1(n535), .A2(n534), .ZN(N836) );
  nd02d1 U497 ( .A1(n533), .A2(n532), .ZN(N835) );
  nd02d1 U498 ( .A1(n531), .A2(n530), .ZN(N834) );
  nd02d1 U499 ( .A1(n529), .A2(n528), .ZN(N833) );
  nd02d1 U500 ( .A1(n527), .A2(n526), .ZN(N832) );
  nd02d1 U501 ( .A1(n525), .A2(n524), .ZN(N831) );
  nd02d1 U502 ( .A1(n523), .A2(n522), .ZN(N830) );
  nd02d1 U503 ( .A1(n521), .A2(n520), .ZN(N829) );
  nd02d1 U504 ( .A1(n519), .A2(n518), .ZN(N828) );
  nd02d1 U505 ( .A1(n517), .A2(n516), .ZN(N827) );
  nd02d1 U506 ( .A1(n515), .A2(n514), .ZN(N826) );
  nd02d1 U507 ( .A1(n513), .A2(n512), .ZN(N825) );
  nd02d1 U508 ( .A1(n511), .A2(n510), .ZN(N824) );
  nd02d1 U509 ( .A1(n509), .A2(n508), .ZN(N823) );
  nd02d1 U510 ( .A1(n507), .A2(n506), .ZN(N822) );
  nd02d1 U511 ( .A1(n505), .A2(n504), .ZN(N821) );
  nd02d1 U512 ( .A1(n503), .A2(n502), .ZN(N820) );
  nd02d1 U513 ( .A1(n501), .A2(n500), .ZN(N819) );
  nd02d1 U514 ( .A1(n499), .A2(n498), .ZN(N818) );
  nd02d1 U515 ( .A1(n497), .A2(n496), .ZN(N817) );
  nd02d1 U516 ( .A1(n495), .A2(n494), .ZN(N816) );
  nd02d1 U517 ( .A1(n493), .A2(n492), .ZN(N815) );
  nd02d1 U518 ( .A1(n491), .A2(n490), .ZN(N814) );
  nd02d1 U519 ( .A1(n489), .A2(n488), .ZN(N813) );
  nd02d1 U520 ( .A1(n487), .A2(n486), .ZN(N812) );
  nd02d1 U521 ( .A1(n485), .A2(n484), .ZN(N811) );
  nd02d1 U522 ( .A1(n483), .A2(n482), .ZN(N810) );
  nd02d1 U523 ( .A1(n481), .A2(n480), .ZN(N809) );
  nd02d1 U524 ( .A1(n479), .A2(n478), .ZN(N808) );
  nd02d1 U525 ( .A1(n477), .A2(n476), .ZN(N807) );
  inv0d1 U526 ( .I(wr_addr_1_), .ZN(n471) );
  inv0d1 U527 ( .I(wr_addr_2_), .ZN(n470) );
  inv0d1 U528 ( .I(wr_addr_0_), .ZN(n468) );
  lanlq1 LOCKUP ( .D(data_out_sync_31_), .EN(fifo_clk_pop), .Q(test_so1) );
endmodule


module SDRAM_FIFO_0 ( fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, 
        fifo_push_req_n, fifo_pop_req_n, fifo_data_in, push_empty_fifo, 
        push_ae_fifo, push_hf_fifo, push_af_fifo, push_full_fifo, 
        push_error_fifo, pop_empty_fifo, pop_ae_fifo, pop_hf_fifo, pop_af_fifo, 
        pop_full_fifo, pop_error_fifo, data_out_fifo, test_se, test_si1, 
        test_si2, test_si3, test_si4, test_so1, test_so2, test_so4 );
  input [31:0] fifo_data_in;
  output [31:0] data_out_fifo;
  input fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, fifo_push_req_n,
         fifo_pop_req_n, test_se, test_si1, test_si2, test_si3, test_si4;
  output push_empty_fifo, push_ae_fifo, push_hf_fifo, push_af_fifo,
         push_full_fifo, push_error_fifo, pop_empty_fifo, pop_ae_fifo,
         pop_hf_fifo, pop_af_fifo, pop_full_fifo, pop_error_fifo, test_so1,
         test_so2, test_so4;
  wire   we_n, reg_array_255_, reg_array_254_, reg_array_253_, reg_array_252_,
         reg_array_251_, reg_array_250_, reg_array_249_, reg_array_248_,
         reg_array_247_, reg_array_246_, reg_array_245_, reg_array_244_,
         reg_array_243_, reg_array_242_, reg_array_241_, reg_array_240_,
         reg_array_239_, reg_array_238_, reg_array_237_, reg_array_236_,
         reg_array_235_, reg_array_234_, reg_array_233_, reg_array_232_,
         reg_array_231_, reg_array_230_, reg_array_229_, reg_array_228_,
         reg_array_227_, reg_array_226_, reg_array_225_, reg_array_224_,
         reg_array_223_, reg_array_222_, reg_array_221_, reg_array_220_,
         reg_array_219_, reg_array_218_, reg_array_217_, reg_array_216_,
         reg_array_215_, reg_array_214_, reg_array_213_, reg_array_212_,
         reg_array_211_, reg_array_210_, reg_array_209_, reg_array_208_,
         reg_array_207_, reg_array_206_, reg_array_205_, reg_array_204_,
         reg_array_203_, reg_array_202_, reg_array_201_, reg_array_200_,
         reg_array_199_, reg_array_198_, reg_array_197_, reg_array_196_,
         reg_array_195_, reg_array_194_, reg_array_193_, reg_array_192_,
         reg_array_191_, reg_array_190_, reg_array_189_, reg_array_188_,
         reg_array_187_, reg_array_186_, reg_array_185_, reg_array_184_,
         reg_array_183_, reg_array_182_, reg_array_181_, reg_array_180_,
         reg_array_179_, reg_array_178_, reg_array_177_, reg_array_176_,
         reg_array_175_, reg_array_174_, reg_array_173_, reg_array_172_,
         reg_array_171_, reg_array_170_, reg_array_169_, reg_array_168_,
         reg_array_167_, reg_array_166_, reg_array_165_, reg_array_163_,
         reg_array_162_, reg_array_161_, reg_array_160_, reg_array_159_,
         reg_array_158_, reg_array_157_, reg_array_156_, reg_array_155_,
         reg_array_154_, reg_array_153_, reg_array_152_, reg_array_151_,
         reg_array_150_, reg_array_149_, reg_array_148_, reg_array_147_,
         reg_array_146_, reg_array_145_, reg_array_144_, reg_array_143_,
         reg_array_142_, reg_array_141_, reg_array_140_, reg_array_139_,
         reg_array_138_, reg_array_137_, reg_array_136_, reg_array_135_,
         reg_array_134_, reg_array_133_, reg_array_132_, reg_array_131_,
         reg_array_130_, reg_array_129_, reg_array_128_, reg_array_127_,
         reg_array_126_, reg_array_125_, reg_array_124_, reg_array_123_,
         reg_array_122_, reg_array_121_, reg_array_120_, reg_array_119_,
         reg_array_118_, reg_array_117_, reg_array_116_, reg_array_115_,
         reg_array_114_, reg_array_113_, reg_array_112_, reg_array_111_,
         reg_array_110_, reg_array_109_, reg_array_108_, reg_array_107_,
         reg_array_106_, reg_array_105_, reg_array_104_, reg_array_103_,
         reg_array_102_, reg_array_101_, reg_array_100_, reg_array_99_,
         reg_array_98_, reg_array_97_, reg_array_96_, reg_array_95_,
         reg_array_94_, reg_array_93_, reg_array_92_, reg_array_91_,
         reg_array_90_, reg_array_89_, reg_array_88_, reg_array_87_,
         reg_array_86_, reg_array_85_, reg_array_84_, reg_array_83_,
         reg_array_82_, reg_array_81_, reg_array_80_, reg_array_79_,
         reg_array_78_, reg_array_77_, reg_array_76_, reg_array_75_,
         reg_array_74_, reg_array_73_, reg_array_72_, reg_array_71_,
         reg_array_70_, reg_array_69_, reg_array_68_, reg_array_67_,
         reg_array_66_, reg_array_65_, reg_array_64_, reg_array_63_,
         reg_array_62_, reg_array_61_, reg_array_60_, reg_array_59_,
         reg_array_58_, reg_array_57_, reg_array_56_, reg_array_55_,
         reg_array_54_, reg_array_53_, reg_array_52_, reg_array_51_,
         reg_array_50_, reg_array_49_, reg_array_48_, reg_array_47_,
         reg_array_46_, reg_array_45_, reg_array_44_, reg_array_43_,
         reg_array_42_, reg_array_41_, reg_array_40_, reg_array_39_,
         reg_array_38_, reg_array_37_, reg_array_36_, reg_array_35_,
         reg_array_34_, reg_array_33_, reg_array_32_, reg_array_30_,
         reg_array_29_, reg_array_28_, reg_array_27_, reg_array_26_,
         reg_array_25_, reg_array_24_, reg_array_23_, reg_array_22_,
         reg_array_21_, reg_array_20_, reg_array_19_, reg_array_18_,
         reg_array_17_, reg_array_16_, reg_array_15_, reg_array_14_,
         reg_array_13_, reg_array_12_, reg_array_11_, reg_array_10_,
         reg_array_9_, reg_array_8_, reg_array_7_, reg_array_6_, reg_array_5_,
         reg_array_4_, reg_array_3_, reg_array_2_, reg_array_1_, reg_array_0_,
         N729, N731, N733, N735, N737, N739, N741, N743, N745, N747, N749,
         N751, N753, N755, N757, N759, N761, N763, N765, N767, N769, N771,
         N773, N775, N777, N779, N781, N783, N785, N787, N789, N791, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838,
         data_out_sync_30_, data_out_sync_29_, data_out_sync_28_,
         data_out_sync_27_, data_out_sync_26_, data_out_sync_25_,
         data_out_sync_24_, data_out_sync_23_, data_out_sync_22_,
         data_out_sync_21_, data_out_sync_20_, data_out_sync_19_,
         data_out_sync_18_, data_out_sync_17_, data_out_sync_16_,
         data_out_sync_15_, data_out_sync_14_, data_out_sync_13_,
         data_out_sync_12_, data_out_sync_11_, data_out_sync_10_,
         data_out_sync_9_, data_out_sync_8_, data_out_sync_7_,
         data_out_sync_6_, data_out_sync_5_, data_out_sync_4_,
         data_out_sync_3_, data_out_sync_2_, data_out_sync_1_,
         data_out_sync_0_, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n1,
         n97, n130, n163, n196, n229, n262, n295, n328, n404, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n465, n468, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16;
  wire   [2:0] wr_addr;
  wire   [2:0] rd_addr;

  an03d1 U363 ( .A1(n402), .A2(n403), .A3(rd_addr[2]), .Z(n335) );
  an03d1 U364 ( .A1(rd_addr[0]), .A2(n403), .A3(rd_addr[2]), .Z(n334) );
  an03d1 U365 ( .A1(rd_addr[1]), .A2(n402), .A3(rd_addr[2]), .Z(n333) );
  an03d1 U366 ( .A1(rd_addr[1]), .A2(rd_addr[0]), .A3(rd_addr[2]), .Z(n332) );
  an02d1 U379 ( .A1(fifo_rst_n), .A2(fifo_data_in[31]), .Z(N791) );
  an02d1 U380 ( .A1(fifo_data_in[30]), .A2(fifo_rst_n), .Z(N789) );
  an02d1 U381 ( .A1(fifo_data_in[29]), .A2(fifo_rst_n), .Z(N787) );
  an02d1 U382 ( .A1(fifo_data_in[28]), .A2(fifo_rst_n), .Z(N785) );
  an02d1 U383 ( .A1(fifo_data_in[27]), .A2(fifo_rst_n), .Z(N783) );
  an02d1 U384 ( .A1(fifo_data_in[26]), .A2(fifo_rst_n), .Z(N781) );
  an02d1 U385 ( .A1(fifo_data_in[25]), .A2(fifo_rst_n), .Z(N779) );
  an02d1 U386 ( .A1(fifo_data_in[24]), .A2(fifo_rst_n), .Z(N777) );
  an02d1 U387 ( .A1(fifo_data_in[23]), .A2(fifo_rst_n), .Z(N775) );
  an02d1 U388 ( .A1(fifo_data_in[22]), .A2(fifo_rst_n), .Z(N773) );
  an02d1 U389 ( .A1(fifo_data_in[21]), .A2(fifo_rst_n), .Z(N771) );
  an02d1 U390 ( .A1(fifo_data_in[20]), .A2(fifo_rst_n), .Z(N769) );
  an02d1 U391 ( .A1(fifo_data_in[19]), .A2(fifo_rst_n), .Z(N767) );
  an02d1 U392 ( .A1(fifo_data_in[18]), .A2(fifo_rst_n), .Z(N765) );
  an02d1 U393 ( .A1(fifo_data_in[17]), .A2(fifo_rst_n), .Z(N763) );
  an02d1 U394 ( .A1(fifo_data_in[16]), .A2(fifo_rst_n), .Z(N761) );
  an02d1 U395 ( .A1(fifo_data_in[15]), .A2(fifo_rst_n), .Z(N759) );
  an02d1 U396 ( .A1(fifo_data_in[14]), .A2(fifo_rst_n), .Z(N757) );
  an02d1 U397 ( .A1(fifo_data_in[13]), .A2(fifo_rst_n), .Z(N755) );
  an02d1 U398 ( .A1(fifo_data_in[12]), .A2(fifo_rst_n), .Z(N753) );
  an02d1 U399 ( .A1(fifo_data_in[11]), .A2(fifo_rst_n), .Z(N751) );
  an02d1 U400 ( .A1(fifo_data_in[10]), .A2(fifo_rst_n), .Z(N749) );
  an02d1 U401 ( .A1(fifo_data_in[9]), .A2(fifo_rst_n), .Z(N747) );
  an02d1 U402 ( .A1(fifo_data_in[8]), .A2(fifo_rst_n), .Z(N745) );
  an02d1 U403 ( .A1(fifo_data_in[7]), .A2(fifo_rst_n), .Z(N743) );
  an02d1 U404 ( .A1(fifo_data_in[6]), .A2(fifo_rst_n), .Z(N741) );
  an02d1 U405 ( .A1(fifo_data_in[5]), .A2(fifo_rst_n), .Z(N739) );
  an02d1 U406 ( .A1(fifo_data_in[4]), .A2(fifo_rst_n), .Z(N737) );
  an02d1 U407 ( .A1(fifo_data_in[3]), .A2(fifo_rst_n), .Z(N735) );
  an02d1 U408 ( .A1(fifo_data_in[2]), .A2(fifo_rst_n), .Z(N733) );
  an02d1 U409 ( .A1(fifo_data_in[1]), .A2(fifo_rst_n), .Z(N731) );
  an02d1 U410 ( .A1(fifo_data_in[0]), .A2(fifo_rst_n), .Z(N729) );
  aoi2222d1 U413 ( .A1(reg_array_0_), .A2(n438), .B1(reg_array_32_), .B2(n435), 
        .C1(reg_array_64_), .C2(n432), .D1(reg_array_96_), .D2(n429), .ZN(n331) );
  aoi2222d1 U414 ( .A1(reg_array_128_), .A2(n426), .B1(reg_array_160_), .B2(
        n423), .C1(reg_array_192_), .C2(n420), .D1(reg_array_224_), .D2(n417), 
        .ZN(n330) );
  aoi2222d1 U415 ( .A1(reg_array_1_), .A2(n438), .B1(reg_array_33_), .B2(n435), 
        .C1(reg_array_65_), .C2(n432), .D1(reg_array_97_), .D2(n429), .ZN(n341) );
  aoi2222d1 U416 ( .A1(reg_array_129_), .A2(n426), .B1(reg_array_161_), .B2(
        n423), .C1(reg_array_193_), .C2(n420), .D1(reg_array_225_), .D2(n417), 
        .ZN(n340) );
  aoi2222d1 U417 ( .A1(reg_array_2_), .A2(n438), .B1(reg_array_34_), .B2(n435), 
        .C1(reg_array_66_), .C2(n432), .D1(reg_array_98_), .D2(n429), .ZN(n343) );
  aoi2222d1 U418 ( .A1(reg_array_130_), .A2(n426), .B1(reg_array_162_), .B2(
        n423), .C1(reg_array_194_), .C2(n420), .D1(reg_array_226_), .D2(n417), 
        .ZN(n342) );
  aoi2222d1 U419 ( .A1(reg_array_3_), .A2(n438), .B1(reg_array_35_), .B2(n435), 
        .C1(reg_array_67_), .C2(n432), .D1(reg_array_99_), .D2(n429), .ZN(n345) );
  aoi2222d1 U420 ( .A1(reg_array_131_), .A2(n426), .B1(reg_array_163_), .B2(
        n423), .C1(reg_array_195_), .C2(n420), .D1(reg_array_227_), .D2(n417), 
        .ZN(n344) );
  aoi2222d1 U421 ( .A1(reg_array_4_), .A2(n438), .B1(reg_array_36_), .B2(n435), 
        .C1(reg_array_68_), .C2(n432), .D1(reg_array_100_), .D2(n429), .ZN(
        n347) );
  aoi2222d1 U422 ( .A1(reg_array_132_), .A2(n426), .B1(test_so2), .B2(n423), 
        .C1(reg_array_196_), .C2(n420), .D1(reg_array_228_), .D2(n417), .ZN(
        n346) );
  aoi2222d1 U423 ( .A1(reg_array_5_), .A2(n438), .B1(reg_array_37_), .B2(n435), 
        .C1(reg_array_69_), .C2(n432), .D1(reg_array_101_), .D2(n429), .ZN(
        n349) );
  aoi2222d1 U424 ( .A1(reg_array_133_), .A2(n426), .B1(reg_array_165_), .B2(
        n423), .C1(reg_array_197_), .C2(n420), .D1(reg_array_229_), .D2(n417), 
        .ZN(n348) );
  aoi2222d1 U425 ( .A1(reg_array_6_), .A2(n438), .B1(reg_array_38_), .B2(n435), 
        .C1(reg_array_70_), .C2(n432), .D1(reg_array_102_), .D2(n429), .ZN(
        n351) );
  aoi2222d1 U426 ( .A1(reg_array_134_), .A2(n426), .B1(reg_array_166_), .B2(
        n423), .C1(reg_array_198_), .C2(n420), .D1(reg_array_230_), .D2(n417), 
        .ZN(n350) );
  aoi2222d1 U427 ( .A1(reg_array_7_), .A2(n438), .B1(reg_array_39_), .B2(n435), 
        .C1(reg_array_71_), .C2(n432), .D1(reg_array_103_), .D2(n429), .ZN(
        n353) );
  aoi2222d1 U428 ( .A1(reg_array_135_), .A2(n426), .B1(reg_array_167_), .B2(
        n423), .C1(reg_array_199_), .C2(n420), .D1(reg_array_231_), .D2(n417), 
        .ZN(n352) );
  aoi2222d1 U429 ( .A1(reg_array_8_), .A2(n438), .B1(reg_array_40_), .B2(n435), 
        .C1(reg_array_72_), .C2(n432), .D1(reg_array_104_), .D2(n429), .ZN(
        n355) );
  aoi2222d1 U430 ( .A1(reg_array_136_), .A2(n426), .B1(reg_array_168_), .B2(
        n423), .C1(reg_array_200_), .C2(n420), .D1(reg_array_232_), .D2(n417), 
        .ZN(n354) );
  aoi2222d1 U431 ( .A1(reg_array_9_), .A2(n438), .B1(reg_array_41_), .B2(n435), 
        .C1(reg_array_73_), .C2(n432), .D1(reg_array_105_), .D2(n429), .ZN(
        n357) );
  aoi2222d1 U432 ( .A1(reg_array_137_), .A2(n426), .B1(reg_array_169_), .B2(
        n423), .C1(reg_array_201_), .C2(n420), .D1(reg_array_233_), .D2(n417), 
        .ZN(n356) );
  aoi2222d1 U433 ( .A1(reg_array_10_), .A2(n437), .B1(reg_array_42_), .B2(n434), .C1(reg_array_74_), .C2(n431), .D1(reg_array_106_), .D2(n428), .ZN(n359) );
  aoi2222d1 U434 ( .A1(reg_array_138_), .A2(n425), .B1(reg_array_170_), .B2(
        n422), .C1(reg_array_202_), .C2(n419), .D1(reg_array_234_), .D2(n416), 
        .ZN(n358) );
  aoi2222d1 U435 ( .A1(reg_array_11_), .A2(n437), .B1(reg_array_43_), .B2(n434), .C1(reg_array_75_), .C2(n431), .D1(reg_array_107_), .D2(n428), .ZN(n361) );
  aoi2222d1 U436 ( .A1(reg_array_139_), .A2(n425), .B1(reg_array_171_), .B2(
        n422), .C1(reg_array_203_), .C2(n419), .D1(reg_array_235_), .D2(n416), 
        .ZN(n360) );
  aoi2222d1 U437 ( .A1(reg_array_12_), .A2(n437), .B1(reg_array_44_), .B2(n434), .C1(reg_array_76_), .C2(n431), .D1(reg_array_108_), .D2(n428), .ZN(n363) );
  aoi2222d1 U438 ( .A1(reg_array_140_), .A2(n425), .B1(reg_array_172_), .B2(
        n422), .C1(reg_array_204_), .C2(n419), .D1(reg_array_236_), .D2(n416), 
        .ZN(n362) );
  aoi2222d1 U439 ( .A1(reg_array_13_), .A2(n437), .B1(reg_array_45_), .B2(n434), .C1(reg_array_77_), .C2(n431), .D1(reg_array_109_), .D2(n428), .ZN(n365) );
  aoi2222d1 U440 ( .A1(reg_array_141_), .A2(n425), .B1(reg_array_173_), .B2(
        n422), .C1(reg_array_205_), .C2(n419), .D1(reg_array_237_), .D2(n416), 
        .ZN(n364) );
  aoi2222d1 U441 ( .A1(reg_array_14_), .A2(n437), .B1(reg_array_46_), .B2(n434), .C1(reg_array_78_), .C2(n431), .D1(reg_array_110_), .D2(n428), .ZN(n367) );
  aoi2222d1 U442 ( .A1(reg_array_142_), .A2(n425), .B1(reg_array_174_), .B2(
        n422), .C1(reg_array_206_), .C2(n419), .D1(reg_array_238_), .D2(n416), 
        .ZN(n366) );
  aoi2222d1 U443 ( .A1(reg_array_15_), .A2(n437), .B1(reg_array_47_), .B2(n434), .C1(reg_array_79_), .C2(n431), .D1(reg_array_111_), .D2(n428), .ZN(n369) );
  aoi2222d1 U444 ( .A1(reg_array_143_), .A2(n425), .B1(reg_array_175_), .B2(
        n422), .C1(reg_array_207_), .C2(n419), .D1(reg_array_239_), .D2(n416), 
        .ZN(n368) );
  aoi2222d1 U445 ( .A1(reg_array_16_), .A2(n437), .B1(reg_array_48_), .B2(n434), .C1(reg_array_80_), .C2(n431), .D1(reg_array_112_), .D2(n428), .ZN(n371) );
  aoi2222d1 U446 ( .A1(reg_array_144_), .A2(n425), .B1(reg_array_176_), .B2(
        n422), .C1(reg_array_208_), .C2(n419), .D1(reg_array_240_), .D2(n416), 
        .ZN(n370) );
  aoi2222d1 U447 ( .A1(reg_array_17_), .A2(n437), .B1(reg_array_49_), .B2(n434), .C1(reg_array_81_), .C2(n431), .D1(reg_array_113_), .D2(n428), .ZN(n373) );
  aoi2222d1 U448 ( .A1(reg_array_145_), .A2(n425), .B1(reg_array_177_), .B2(
        n422), .C1(reg_array_209_), .C2(n419), .D1(reg_array_241_), .D2(n416), 
        .ZN(n372) );
  aoi2222d1 U449 ( .A1(reg_array_18_), .A2(n437), .B1(reg_array_50_), .B2(n434), .C1(reg_array_82_), .C2(n431), .D1(reg_array_114_), .D2(n428), .ZN(n375) );
  aoi2222d1 U450 ( .A1(reg_array_146_), .A2(n425), .B1(reg_array_178_), .B2(
        n422), .C1(reg_array_210_), .C2(n419), .D1(reg_array_242_), .D2(n416), 
        .ZN(n374) );
  aoi2222d1 U451 ( .A1(reg_array_19_), .A2(n437), .B1(reg_array_51_), .B2(n434), .C1(reg_array_83_), .C2(n431), .D1(reg_array_115_), .D2(n428), .ZN(n377) );
  aoi2222d1 U452 ( .A1(reg_array_147_), .A2(n425), .B1(reg_array_179_), .B2(
        n422), .C1(reg_array_211_), .C2(n419), .D1(reg_array_243_), .D2(n416), 
        .ZN(n376) );
  aoi2222d1 U453 ( .A1(reg_array_20_), .A2(n437), .B1(reg_array_52_), .B2(n434), .C1(reg_array_84_), .C2(n431), .D1(reg_array_116_), .D2(n428), .ZN(n379) );
  aoi2222d1 U454 ( .A1(reg_array_148_), .A2(n425), .B1(reg_array_180_), .B2(
        n422), .C1(reg_array_212_), .C2(n419), .D1(reg_array_244_), .D2(n416), 
        .ZN(n378) );
  aoi2222d1 U455 ( .A1(reg_array_21_), .A2(n436), .B1(reg_array_53_), .B2(n433), .C1(reg_array_85_), .C2(n430), .D1(reg_array_117_), .D2(n427), .ZN(n381) );
  aoi2222d1 U456 ( .A1(reg_array_149_), .A2(n424), .B1(reg_array_181_), .B2(
        n421), .C1(reg_array_213_), .C2(n418), .D1(reg_array_245_), .D2(n404), 
        .ZN(n380) );
  aoi2222d1 U457 ( .A1(reg_array_22_), .A2(n436), .B1(reg_array_54_), .B2(n433), .C1(reg_array_86_), .C2(n430), .D1(reg_array_118_), .D2(n427), .ZN(n383) );
  aoi2222d1 U458 ( .A1(reg_array_150_), .A2(n424), .B1(reg_array_182_), .B2(
        n421), .C1(reg_array_214_), .C2(n418), .D1(reg_array_246_), .D2(n404), 
        .ZN(n382) );
  aoi2222d1 U459 ( .A1(reg_array_23_), .A2(n436), .B1(reg_array_55_), .B2(n433), .C1(reg_array_87_), .C2(n430), .D1(reg_array_119_), .D2(n427), .ZN(n385) );
  aoi2222d1 U460 ( .A1(reg_array_151_), .A2(n424), .B1(reg_array_183_), .B2(
        n421), .C1(reg_array_215_), .C2(n418), .D1(reg_array_247_), .D2(n404), 
        .ZN(n384) );
  aoi2222d1 U461 ( .A1(reg_array_24_), .A2(n436), .B1(reg_array_56_), .B2(n433), .C1(reg_array_88_), .C2(n430), .D1(reg_array_120_), .D2(n427), .ZN(n387) );
  aoi2222d1 U462 ( .A1(reg_array_152_), .A2(n424), .B1(reg_array_184_), .B2(
        n421), .C1(reg_array_216_), .C2(n418), .D1(reg_array_248_), .D2(n404), 
        .ZN(n386) );
  aoi2222d1 U463 ( .A1(reg_array_25_), .A2(n436), .B1(reg_array_57_), .B2(n433), .C1(reg_array_89_), .C2(n430), .D1(reg_array_121_), .D2(n427), .ZN(n389) );
  aoi2222d1 U464 ( .A1(reg_array_153_), .A2(n424), .B1(reg_array_185_), .B2(
        n421), .C1(reg_array_217_), .C2(n418), .D1(reg_array_249_), .D2(n404), 
        .ZN(n388) );
  aoi2222d1 U465 ( .A1(reg_array_26_), .A2(n436), .B1(reg_array_58_), .B2(n433), .C1(reg_array_90_), .C2(n430), .D1(reg_array_122_), .D2(n427), .ZN(n391) );
  aoi2222d1 U466 ( .A1(reg_array_154_), .A2(n424), .B1(reg_array_186_), .B2(
        n421), .C1(reg_array_218_), .C2(n418), .D1(reg_array_250_), .D2(n404), 
        .ZN(n390) );
  aoi2222d1 U467 ( .A1(reg_array_27_), .A2(n436), .B1(reg_array_59_), .B2(n433), .C1(reg_array_91_), .C2(n430), .D1(reg_array_123_), .D2(n427), .ZN(n393) );
  aoi2222d1 U468 ( .A1(reg_array_155_), .A2(n424), .B1(reg_array_187_), .B2(
        n421), .C1(reg_array_219_), .C2(n418), .D1(reg_array_251_), .D2(n404), 
        .ZN(n392) );
  aoi2222d1 U469 ( .A1(reg_array_28_), .A2(n436), .B1(reg_array_60_), .B2(n433), .C1(reg_array_92_), .C2(n430), .D1(reg_array_124_), .D2(n427), .ZN(n395) );
  aoi2222d1 U470 ( .A1(reg_array_156_), .A2(n424), .B1(reg_array_188_), .B2(
        n421), .C1(reg_array_220_), .C2(n418), .D1(reg_array_252_), .D2(n404), 
        .ZN(n394) );
  aoi2222d1 U471 ( .A1(reg_array_29_), .A2(n436), .B1(reg_array_61_), .B2(n433), .C1(reg_array_93_), .C2(n430), .D1(reg_array_125_), .D2(n427), .ZN(n397) );
  aoi2222d1 U472 ( .A1(reg_array_157_), .A2(n424), .B1(reg_array_189_), .B2(
        n421), .C1(reg_array_221_), .C2(n418), .D1(reg_array_253_), .D2(n404), 
        .ZN(n396) );
  aoi2222d1 U473 ( .A1(reg_array_30_), .A2(n436), .B1(reg_array_62_), .B2(n433), .C1(reg_array_94_), .C2(n430), .D1(reg_array_126_), .D2(n427), .ZN(n399) );
  aoi2222d1 U474 ( .A1(reg_array_158_), .A2(n424), .B1(reg_array_190_), .B2(
        n421), .C1(reg_array_222_), .C2(n418), .D1(reg_array_254_), .D2(n404), 
        .ZN(n398) );
  aoi2222d1 U475 ( .A1(test_so4), .A2(n436), .B1(reg_array_63_), .B2(n433), 
        .C1(reg_array_95_), .C2(n430), .D1(reg_array_127_), .D2(n427), .ZN(
        n401) );
  aoi2222d1 U476 ( .A1(reg_array_159_), .A2(n424), .B1(reg_array_191_), .B2(
        n421), .C1(reg_array_223_), .C2(n418), .D1(reg_array_255_), .D2(n404), 
        .ZN(n400) );
  nr03d0 U477 ( .A1(rd_addr[1]), .A2(rd_addr[2]), .A3(rd_addr[0]), .ZN(n339)
         );
  nr03d0 U478 ( .A1(rd_addr[1]), .A2(rd_addr[2]), .A3(n402), .ZN(n338) );
  nr03d0 U479 ( .A1(rd_addr[0]), .A2(rd_addr[2]), .A3(n403), .ZN(n337) );
  nr03d0 U480 ( .A1(n402), .A2(rd_addr[2]), .A3(n403), .ZN(n336) );
  nd04d0 U482 ( .A1(wr_addr[0]), .A2(n406), .A3(n407), .A4(n408), .ZN(n405) );
  nd04d0 U483 ( .A1(wr_addr[1]), .A2(n406), .A3(n410), .A4(n408), .ZN(n409) );
  nd04d0 U484 ( .A1(wr_addr[1]), .A2(wr_addr[0]), .A3(n406), .A4(n408), .ZN(
        n411) );
  nd04d0 U485 ( .A1(wr_addr[2]), .A2(n406), .A3(n410), .A4(n407), .ZN(n412) );
  nd04d0 U486 ( .A1(wr_addr[2]), .A2(wr_addr[0]), .A3(n406), .A4(n407), .ZN(
        n413) );
  nd04d0 U487 ( .A1(wr_addr[2]), .A2(wr_addr[1]), .A3(n406), .A4(n410), .ZN(
        n414) );
  nd04d0 U488 ( .A1(wr_addr[2]), .A2(wr_addr[1]), .A3(wr_addr[0]), .A4(n406), 
        .ZN(n415) );
  SDRAM_FIFO_0_DW_fifoctl_s2_sf_0 SD_FIFO_CTL ( .clk_push(fifo_clk_push), 
        .clk_pop(fifo_clk_pop), .rst_n(fifo_rst_n), .push_req_n(
        fifo_push_req_n), .pop_req_n(fifo_pop_req_n), .we_n(we_n), 
        .push_empty(push_empty_fifo), .push_ae(push_ae_fifo), .push_hf(
        push_hf_fifo), .push_af(push_af_fifo), .push_full(push_full_fifo), 
        .push_error(push_error_fifo), .pop_empty(pop_empty_fifo), .pop_ae(
        pop_ae_fifo), .pop_hf(pop_hf_fifo), .pop_af(pop_af_fifo), .pop_full(
        pop_full_fifo), .pop_error(pop_error_fifo), .wr_addr(wr_addr), 
        .rd_addr(rd_addr), .push_word_count({SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12}), .pop_word_count({SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16}), .test(test_mode), .test_si1(test_si2), 
        .test_si2(test_si3), .test_se(test_se), .test_so1(n468), .test_so2(
        n465) );
  senrq1 reg_array_reg_0__31_ ( .D(N791), .SD(reg_array_254_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_255_) );
  senrq1 reg_array_reg_0__30_ ( .D(N789), .SD(reg_array_253_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_254_) );
  senrq1 reg_array_reg_0__29_ ( .D(N787), .SD(reg_array_252_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_253_) );
  senrq1 reg_array_reg_0__28_ ( .D(N785), .SD(reg_array_251_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_252_) );
  senrq1 reg_array_reg_0__27_ ( .D(N783), .SD(reg_array_250_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_251_) );
  senrq1 reg_array_reg_0__26_ ( .D(N781), .SD(reg_array_249_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_250_) );
  senrq1 reg_array_reg_0__25_ ( .D(N779), .SD(reg_array_248_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_249_) );
  senrq1 reg_array_reg_0__24_ ( .D(N777), .SD(reg_array_247_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_248_) );
  senrq1 reg_array_reg_0__23_ ( .D(N775), .SD(reg_array_246_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_247_) );
  senrq1 reg_array_reg_0__22_ ( .D(N773), .SD(reg_array_245_), .ENN(n441), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_246_) );
  senrq1 reg_array_reg_0__21_ ( .D(N771), .SD(reg_array_244_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_245_) );
  senrq1 reg_array_reg_0__20_ ( .D(N769), .SD(reg_array_243_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_244_) );
  senrq1 reg_array_reg_0__19_ ( .D(N767), .SD(reg_array_242_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_243_) );
  senrq1 reg_array_reg_0__18_ ( .D(N765), .SD(reg_array_241_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_242_) );
  senrq1 reg_array_reg_0__17_ ( .D(N763), .SD(reg_array_240_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_241_) );
  senrq1 reg_array_reg_0__16_ ( .D(N761), .SD(reg_array_239_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_240_) );
  senrq1 reg_array_reg_0__15_ ( .D(N759), .SD(reg_array_238_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_239_) );
  senrq1 reg_array_reg_0__14_ ( .D(N757), .SD(reg_array_237_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_238_) );
  senrq1 reg_array_reg_0__13_ ( .D(N755), .SD(reg_array_236_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_237_) );
  senrq1 reg_array_reg_0__12_ ( .D(N753), .SD(reg_array_235_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_236_) );
  senrq1 reg_array_reg_0__11_ ( .D(N751), .SD(reg_array_234_), .ENN(n440), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_235_) );
  senrq1 reg_array_reg_0__10_ ( .D(N749), .SD(reg_array_233_), .ENN(n439), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_234_) );
  senrq1 reg_array_reg_0__9_ ( .D(N747), .SD(reg_array_232_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_233_) );
  senrq1 reg_array_reg_0__8_ ( .D(N745), .SD(reg_array_231_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_232_) );
  senrq1 reg_array_reg_0__7_ ( .D(N743), .SD(reg_array_230_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_231_) );
  senrq1 reg_array_reg_0__6_ ( .D(N741), .SD(reg_array_229_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_230_) );
  senrq1 reg_array_reg_0__5_ ( .D(N739), .SD(reg_array_228_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_229_) );
  senrq1 reg_array_reg_0__4_ ( .D(N737), .SD(reg_array_227_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_228_) );
  senrq1 reg_array_reg_0__3_ ( .D(N735), .SD(reg_array_226_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_227_) );
  senrq1 reg_array_reg_0__2_ ( .D(N733), .SD(reg_array_225_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_226_) );
  senrq1 reg_array_reg_0__1_ ( .D(N731), .SD(reg_array_224_), .ENN(n439), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_225_) );
  senrq1 reg_array_reg_0__0_ ( .D(N729), .SD(n468), .ENN(n439), .SC(test_se), 
        .CP(fifo_clk_push), .Q(reg_array_224_) );
  senrq1 reg_array_reg_1__31_ ( .D(N791), .SD(reg_array_222_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_223_) );
  senrq1 reg_array_reg_1__30_ ( .D(N789), .SD(reg_array_221_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_222_) );
  senrq1 reg_array_reg_1__29_ ( .D(N787), .SD(reg_array_220_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_221_) );
  senrq1 reg_array_reg_1__28_ ( .D(N785), .SD(reg_array_219_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_220_) );
  senrq1 reg_array_reg_1__27_ ( .D(N783), .SD(reg_array_218_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_219_) );
  senrq1 reg_array_reg_1__26_ ( .D(N781), .SD(reg_array_217_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_218_) );
  senrq1 reg_array_reg_1__25_ ( .D(N779), .SD(reg_array_216_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_217_) );
  senrq1 reg_array_reg_1__24_ ( .D(N777), .SD(reg_array_215_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_216_) );
  senrq1 reg_array_reg_1__23_ ( .D(N775), .SD(reg_array_214_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_215_) );
  senrq1 reg_array_reg_1__22_ ( .D(N773), .SD(reg_array_213_), .ENN(n444), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_214_) );
  senrq1 reg_array_reg_1__21_ ( .D(N771), .SD(reg_array_212_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_213_) );
  senrq1 reg_array_reg_1__20_ ( .D(N769), .SD(reg_array_211_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_212_) );
  senrq1 reg_array_reg_1__19_ ( .D(N767), .SD(reg_array_210_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_211_) );
  senrq1 reg_array_reg_1__18_ ( .D(N765), .SD(reg_array_209_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_210_) );
  senrq1 reg_array_reg_1__17_ ( .D(N763), .SD(reg_array_208_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_209_) );
  senrq1 reg_array_reg_1__16_ ( .D(N761), .SD(reg_array_207_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_208_) );
  senrq1 reg_array_reg_1__15_ ( .D(N759), .SD(reg_array_206_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_207_) );
  senrq1 reg_array_reg_1__14_ ( .D(N757), .SD(reg_array_205_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_206_) );
  senrq1 reg_array_reg_1__13_ ( .D(N755), .SD(reg_array_204_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_205_) );
  senrq1 reg_array_reg_1__12_ ( .D(N753), .SD(reg_array_203_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_204_) );
  senrq1 reg_array_reg_1__11_ ( .D(N751), .SD(reg_array_202_), .ENN(n443), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_203_) );
  senrq1 reg_array_reg_1__10_ ( .D(N749), .SD(reg_array_201_), .ENN(n442), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_202_) );
  senrq1 reg_array_reg_1__9_ ( .D(N747), .SD(reg_array_200_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_201_) );
  senrq1 reg_array_reg_1__8_ ( .D(N745), .SD(reg_array_199_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_200_) );
  senrq1 reg_array_reg_1__7_ ( .D(N743), .SD(reg_array_198_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_199_) );
  senrq1 reg_array_reg_1__6_ ( .D(N741), .SD(reg_array_197_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_198_) );
  senrq1 reg_array_reg_1__5_ ( .D(N739), .SD(reg_array_196_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_197_) );
  senrq1 reg_array_reg_1__4_ ( .D(N737), .SD(reg_array_195_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_196_) );
  senrq1 reg_array_reg_1__3_ ( .D(N735), .SD(reg_array_194_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_195_) );
  senrq1 reg_array_reg_1__2_ ( .D(N733), .SD(reg_array_193_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_194_) );
  senrq1 reg_array_reg_1__1_ ( .D(N731), .SD(reg_array_192_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_193_) );
  senrq1 reg_array_reg_1__0_ ( .D(N729), .SD(reg_array_255_), .ENN(n442), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_192_) );
  senrq1 reg_array_reg_2__31_ ( .D(N791), .SD(reg_array_190_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_191_) );
  senrq1 reg_array_reg_2__30_ ( .D(N789), .SD(reg_array_189_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_190_) );
  senrq1 reg_array_reg_2__29_ ( .D(N787), .SD(reg_array_188_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_189_) );
  senrq1 reg_array_reg_2__28_ ( .D(N785), .SD(reg_array_187_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_188_) );
  senrq1 reg_array_reg_2__27_ ( .D(N783), .SD(reg_array_186_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_187_) );
  senrq1 reg_array_reg_2__26_ ( .D(N781), .SD(reg_array_185_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_186_) );
  senrq1 reg_array_reg_2__25_ ( .D(N779), .SD(reg_array_184_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_185_) );
  senrq1 reg_array_reg_2__24_ ( .D(N777), .SD(reg_array_183_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_184_) );
  senrq1 reg_array_reg_2__23_ ( .D(N775), .SD(reg_array_182_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_183_) );
  senrq1 reg_array_reg_2__22_ ( .D(N773), .SD(reg_array_181_), .ENN(n447), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_182_) );
  senrq1 reg_array_reg_2__21_ ( .D(N771), .SD(reg_array_180_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_181_) );
  senrq1 reg_array_reg_2__20_ ( .D(N769), .SD(reg_array_179_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_180_) );
  senrq1 reg_array_reg_2__19_ ( .D(N767), .SD(reg_array_178_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_179_) );
  senrq1 reg_array_reg_2__18_ ( .D(N765), .SD(reg_array_177_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_178_) );
  senrq1 reg_array_reg_2__17_ ( .D(N763), .SD(reg_array_176_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_177_) );
  senrq1 reg_array_reg_2__16_ ( .D(N761), .SD(reg_array_175_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_176_) );
  senrq1 reg_array_reg_2__15_ ( .D(N759), .SD(reg_array_174_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_175_) );
  senrq1 reg_array_reg_2__14_ ( .D(N757), .SD(reg_array_173_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_174_) );
  senrq1 reg_array_reg_2__13_ ( .D(N755), .SD(reg_array_172_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_173_) );
  senrq1 reg_array_reg_2__12_ ( .D(N753), .SD(reg_array_171_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_172_) );
  senrq1 reg_array_reg_2__11_ ( .D(N751), .SD(reg_array_170_), .ENN(n446), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_171_) );
  senrq1 reg_array_reg_2__10_ ( .D(N749), .SD(reg_array_169_), .ENN(n445), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_170_) );
  senrq1 reg_array_reg_2__9_ ( .D(N747), .SD(reg_array_168_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_169_) );
  senrq1 reg_array_reg_2__8_ ( .D(N745), .SD(reg_array_167_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_168_) );
  senrq1 reg_array_reg_2__7_ ( .D(N743), .SD(reg_array_166_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_167_) );
  senrq1 reg_array_reg_2__6_ ( .D(N741), .SD(reg_array_165_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_166_) );
  senrq1 reg_array_reg_2__5_ ( .D(N739), .SD(test_si4), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_165_) );
  senrq1 reg_array_reg_2__4_ ( .D(N737), .SD(reg_array_163_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(test_so2) );
  senrq1 reg_array_reg_2__3_ ( .D(N735), .SD(reg_array_162_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_163_) );
  senrq1 reg_array_reg_2__2_ ( .D(N733), .SD(reg_array_161_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_162_) );
  senrq1 reg_array_reg_2__1_ ( .D(N731), .SD(reg_array_160_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_161_) );
  senrq1 reg_array_reg_2__0_ ( .D(N729), .SD(reg_array_223_), .ENN(n445), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_160_) );
  senrq1 reg_array_reg_3__31_ ( .D(N791), .SD(reg_array_158_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_159_) );
  senrq1 reg_array_reg_3__30_ ( .D(N789), .SD(reg_array_157_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_158_) );
  senrq1 reg_array_reg_3__29_ ( .D(N787), .SD(reg_array_156_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_157_) );
  senrq1 reg_array_reg_3__28_ ( .D(N785), .SD(reg_array_155_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_156_) );
  senrq1 reg_array_reg_3__27_ ( .D(N783), .SD(reg_array_154_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_155_) );
  senrq1 reg_array_reg_3__26_ ( .D(N781), .SD(reg_array_153_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_154_) );
  senrq1 reg_array_reg_3__25_ ( .D(N779), .SD(reg_array_152_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_153_) );
  senrq1 reg_array_reg_3__24_ ( .D(N777), .SD(reg_array_151_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_152_) );
  senrq1 reg_array_reg_3__23_ ( .D(N775), .SD(reg_array_150_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_151_) );
  senrq1 reg_array_reg_3__22_ ( .D(N773), .SD(reg_array_149_), .ENN(n450), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_150_) );
  senrq1 reg_array_reg_3__21_ ( .D(N771), .SD(reg_array_148_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_149_) );
  senrq1 reg_array_reg_3__20_ ( .D(N769), .SD(reg_array_147_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_148_) );
  senrq1 reg_array_reg_3__19_ ( .D(N767), .SD(reg_array_146_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_147_) );
  senrq1 reg_array_reg_3__18_ ( .D(N765), .SD(reg_array_145_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_146_) );
  senrq1 reg_array_reg_3__17_ ( .D(N763), .SD(reg_array_144_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_145_) );
  senrq1 reg_array_reg_3__16_ ( .D(N761), .SD(reg_array_143_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_144_) );
  senrq1 reg_array_reg_3__15_ ( .D(N759), .SD(reg_array_142_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_143_) );
  senrq1 reg_array_reg_3__14_ ( .D(N757), .SD(reg_array_141_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_142_) );
  senrq1 reg_array_reg_3__13_ ( .D(N755), .SD(reg_array_140_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_141_) );
  senrq1 reg_array_reg_3__12_ ( .D(N753), .SD(reg_array_139_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_140_) );
  senrq1 reg_array_reg_3__11_ ( .D(N751), .SD(reg_array_138_), .ENN(n449), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_139_) );
  senrq1 reg_array_reg_3__10_ ( .D(N749), .SD(reg_array_137_), .ENN(n448), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_138_) );
  senrq1 reg_array_reg_3__9_ ( .D(N747), .SD(reg_array_136_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_137_) );
  senrq1 reg_array_reg_3__8_ ( .D(N745), .SD(reg_array_135_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_136_) );
  senrq1 reg_array_reg_3__7_ ( .D(N743), .SD(reg_array_134_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_135_) );
  senrq1 reg_array_reg_3__6_ ( .D(N741), .SD(reg_array_133_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_134_) );
  senrq1 reg_array_reg_3__5_ ( .D(N739), .SD(reg_array_132_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_133_) );
  senrq1 reg_array_reg_3__4_ ( .D(N737), .SD(reg_array_131_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_132_) );
  senrq1 reg_array_reg_3__3_ ( .D(N735), .SD(reg_array_130_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_131_) );
  senrq1 reg_array_reg_3__2_ ( .D(N733), .SD(reg_array_129_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_130_) );
  senrq1 reg_array_reg_3__1_ ( .D(N731), .SD(reg_array_128_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_129_) );
  senrq1 reg_array_reg_3__0_ ( .D(N729), .SD(reg_array_191_), .ENN(n448), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_128_) );
  senrq1 reg_array_reg_4__31_ ( .D(N791), .SD(reg_array_126_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_127_) );
  senrq1 reg_array_reg_4__30_ ( .D(N789), .SD(reg_array_125_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_126_) );
  senrq1 reg_array_reg_4__29_ ( .D(N787), .SD(reg_array_124_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_125_) );
  senrq1 reg_array_reg_4__28_ ( .D(N785), .SD(reg_array_123_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_124_) );
  senrq1 reg_array_reg_4__27_ ( .D(N783), .SD(reg_array_122_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_123_) );
  senrq1 reg_array_reg_4__26_ ( .D(N781), .SD(reg_array_121_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_122_) );
  senrq1 reg_array_reg_4__25_ ( .D(N779), .SD(reg_array_120_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_121_) );
  senrq1 reg_array_reg_4__24_ ( .D(N777), .SD(reg_array_119_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_120_) );
  senrq1 reg_array_reg_4__23_ ( .D(N775), .SD(reg_array_118_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_119_) );
  senrq1 reg_array_reg_4__22_ ( .D(N773), .SD(reg_array_117_), .ENN(n453), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_118_) );
  senrq1 reg_array_reg_4__21_ ( .D(N771), .SD(reg_array_116_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_117_) );
  senrq1 reg_array_reg_4__20_ ( .D(N769), .SD(reg_array_115_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_116_) );
  senrq1 reg_array_reg_4__19_ ( .D(N767), .SD(reg_array_114_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_115_) );
  senrq1 reg_array_reg_4__18_ ( .D(N765), .SD(reg_array_113_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_114_) );
  senrq1 reg_array_reg_4__17_ ( .D(N763), .SD(reg_array_112_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_113_) );
  senrq1 reg_array_reg_4__16_ ( .D(N761), .SD(reg_array_111_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_112_) );
  senrq1 reg_array_reg_4__15_ ( .D(N759), .SD(reg_array_110_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_111_) );
  senrq1 reg_array_reg_4__14_ ( .D(N757), .SD(reg_array_109_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_110_) );
  senrq1 reg_array_reg_4__13_ ( .D(N755), .SD(reg_array_108_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_109_) );
  senrq1 reg_array_reg_4__12_ ( .D(N753), .SD(reg_array_107_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_108_) );
  senrq1 reg_array_reg_4__11_ ( .D(N751), .SD(reg_array_106_), .ENN(n452), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_107_) );
  senrq1 reg_array_reg_4__10_ ( .D(N749), .SD(reg_array_105_), .ENN(n451), 
        .SC(test_se), .CP(fifo_clk_push), .Q(reg_array_106_) );
  senrq1 reg_array_reg_4__9_ ( .D(N747), .SD(reg_array_104_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_105_) );
  senrq1 reg_array_reg_4__8_ ( .D(N745), .SD(reg_array_103_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_104_) );
  senrq1 reg_array_reg_4__7_ ( .D(N743), .SD(reg_array_102_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_103_) );
  senrq1 reg_array_reg_4__6_ ( .D(N741), .SD(reg_array_101_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_102_) );
  senrq1 reg_array_reg_4__5_ ( .D(N739), .SD(reg_array_100_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_101_) );
  senrq1 reg_array_reg_4__4_ ( .D(N737), .SD(reg_array_99_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_100_) );
  senrq1 reg_array_reg_4__3_ ( .D(N735), .SD(reg_array_98_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_99_) );
  senrq1 reg_array_reg_4__2_ ( .D(N733), .SD(reg_array_97_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_98_) );
  senrq1 reg_array_reg_4__1_ ( .D(N731), .SD(reg_array_96_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_97_) );
  senrq1 reg_array_reg_4__0_ ( .D(N729), .SD(reg_array_159_), .ENN(n451), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_96_) );
  senrq1 reg_array_reg_5__31_ ( .D(N791), .SD(reg_array_94_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_95_) );
  senrq1 reg_array_reg_5__30_ ( .D(N789), .SD(reg_array_93_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_94_) );
  senrq1 reg_array_reg_5__29_ ( .D(N787), .SD(reg_array_92_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_93_) );
  senrq1 reg_array_reg_5__28_ ( .D(N785), .SD(reg_array_91_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_92_) );
  senrq1 reg_array_reg_5__27_ ( .D(N783), .SD(reg_array_90_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_91_) );
  senrq1 reg_array_reg_5__26_ ( .D(N781), .SD(reg_array_89_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_90_) );
  senrq1 reg_array_reg_5__25_ ( .D(N779), .SD(reg_array_88_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_89_) );
  senrq1 reg_array_reg_5__24_ ( .D(N777), .SD(reg_array_87_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_88_) );
  senrq1 reg_array_reg_5__23_ ( .D(N775), .SD(reg_array_86_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_87_) );
  senrq1 reg_array_reg_5__22_ ( .D(N773), .SD(reg_array_85_), .ENN(n456), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_86_) );
  senrq1 reg_array_reg_5__21_ ( .D(N771), .SD(reg_array_84_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_85_) );
  senrq1 reg_array_reg_5__20_ ( .D(N769), .SD(reg_array_83_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_84_) );
  senrq1 reg_array_reg_5__19_ ( .D(N767), .SD(reg_array_82_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_83_) );
  senrq1 reg_array_reg_5__18_ ( .D(N765), .SD(reg_array_81_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_82_) );
  senrq1 reg_array_reg_5__17_ ( .D(N763), .SD(reg_array_80_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_81_) );
  senrq1 reg_array_reg_5__16_ ( .D(N761), .SD(reg_array_79_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_80_) );
  senrq1 reg_array_reg_5__15_ ( .D(N759), .SD(reg_array_78_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_79_) );
  senrq1 reg_array_reg_5__14_ ( .D(N757), .SD(reg_array_77_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_78_) );
  senrq1 reg_array_reg_5__13_ ( .D(N755), .SD(reg_array_76_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_77_) );
  senrq1 reg_array_reg_5__12_ ( .D(N753), .SD(reg_array_75_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_76_) );
  senrq1 reg_array_reg_5__11_ ( .D(N751), .SD(reg_array_74_), .ENN(n455), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_75_) );
  senrq1 reg_array_reg_5__10_ ( .D(N749), .SD(reg_array_73_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_74_) );
  senrq1 reg_array_reg_5__9_ ( .D(N747), .SD(reg_array_72_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_73_) );
  senrq1 reg_array_reg_5__8_ ( .D(N745), .SD(reg_array_71_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_72_) );
  senrq1 reg_array_reg_5__7_ ( .D(N743), .SD(reg_array_70_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_71_) );
  senrq1 reg_array_reg_5__6_ ( .D(N741), .SD(reg_array_69_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_70_) );
  senrq1 reg_array_reg_5__5_ ( .D(N739), .SD(reg_array_68_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_69_) );
  senrq1 reg_array_reg_5__4_ ( .D(N737), .SD(reg_array_67_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_68_) );
  senrq1 reg_array_reg_5__3_ ( .D(N735), .SD(reg_array_66_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_67_) );
  senrq1 reg_array_reg_5__2_ ( .D(N733), .SD(reg_array_65_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_66_) );
  senrq1 reg_array_reg_5__1_ ( .D(N731), .SD(reg_array_64_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_65_) );
  senrq1 reg_array_reg_5__0_ ( .D(N729), .SD(reg_array_127_), .ENN(n454), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_64_) );
  senrq1 reg_array_reg_6__31_ ( .D(N791), .SD(reg_array_62_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_63_) );
  senrq1 reg_array_reg_6__30_ ( .D(N789), .SD(reg_array_61_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_62_) );
  senrq1 reg_array_reg_6__29_ ( .D(N787), .SD(reg_array_60_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_61_) );
  senrq1 reg_array_reg_6__28_ ( .D(N785), .SD(reg_array_59_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_60_) );
  senrq1 reg_array_reg_6__27_ ( .D(N783), .SD(reg_array_58_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_59_) );
  senrq1 reg_array_reg_6__26_ ( .D(N781), .SD(reg_array_57_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_58_) );
  senrq1 reg_array_reg_6__25_ ( .D(N779), .SD(reg_array_56_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_57_) );
  senrq1 reg_array_reg_6__24_ ( .D(N777), .SD(reg_array_55_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_56_) );
  senrq1 reg_array_reg_6__23_ ( .D(N775), .SD(reg_array_54_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_55_) );
  senrq1 reg_array_reg_6__22_ ( .D(N773), .SD(reg_array_53_), .ENN(n459), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_54_) );
  senrq1 reg_array_reg_6__21_ ( .D(N771), .SD(reg_array_52_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_53_) );
  senrq1 reg_array_reg_6__20_ ( .D(N769), .SD(reg_array_51_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_52_) );
  senrq1 reg_array_reg_6__19_ ( .D(N767), .SD(reg_array_50_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_51_) );
  senrq1 reg_array_reg_6__18_ ( .D(N765), .SD(reg_array_49_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_50_) );
  senrq1 reg_array_reg_6__17_ ( .D(N763), .SD(reg_array_48_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_49_) );
  senrq1 reg_array_reg_6__16_ ( .D(N761), .SD(reg_array_47_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_48_) );
  senrq1 reg_array_reg_6__15_ ( .D(N759), .SD(reg_array_46_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_47_) );
  senrq1 reg_array_reg_6__14_ ( .D(N757), .SD(reg_array_45_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_46_) );
  senrq1 reg_array_reg_6__13_ ( .D(N755), .SD(reg_array_44_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_45_) );
  senrq1 reg_array_reg_6__12_ ( .D(N753), .SD(reg_array_43_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_44_) );
  senrq1 reg_array_reg_6__11_ ( .D(N751), .SD(reg_array_42_), .ENN(n458), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_43_) );
  senrq1 reg_array_reg_6__10_ ( .D(N749), .SD(reg_array_41_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_42_) );
  senrq1 reg_array_reg_6__9_ ( .D(N747), .SD(reg_array_40_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_41_) );
  senrq1 reg_array_reg_6__8_ ( .D(N745), .SD(reg_array_39_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_40_) );
  senrq1 reg_array_reg_6__7_ ( .D(N743), .SD(reg_array_38_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_39_) );
  senrq1 reg_array_reg_6__6_ ( .D(N741), .SD(reg_array_37_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_38_) );
  senrq1 reg_array_reg_6__5_ ( .D(N739), .SD(reg_array_36_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_37_) );
  senrq1 reg_array_reg_6__4_ ( .D(N737), .SD(reg_array_35_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_36_) );
  senrq1 reg_array_reg_6__3_ ( .D(N735), .SD(reg_array_34_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_35_) );
  senrq1 reg_array_reg_6__2_ ( .D(N733), .SD(reg_array_33_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_34_) );
  senrq1 reg_array_reg_6__1_ ( .D(N731), .SD(reg_array_32_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_33_) );
  senrq1 reg_array_reg_6__0_ ( .D(N729), .SD(reg_array_95_), .ENN(n457), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_32_) );
  senrq1 reg_array_reg_7__31_ ( .D(N791), .SD(reg_array_30_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(test_so4) );
  senrq1 reg_array_reg_7__30_ ( .D(N789), .SD(reg_array_29_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_30_) );
  senrq1 reg_array_reg_7__29_ ( .D(N787), .SD(reg_array_28_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_29_) );
  senrq1 reg_array_reg_7__28_ ( .D(N785), .SD(reg_array_27_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_28_) );
  senrq1 reg_array_reg_7__27_ ( .D(N783), .SD(reg_array_26_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_27_) );
  senrq1 reg_array_reg_7__26_ ( .D(N781), .SD(reg_array_25_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_26_) );
  senrq1 reg_array_reg_7__25_ ( .D(N779), .SD(reg_array_24_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_25_) );
  senrq1 reg_array_reg_7__24_ ( .D(N777), .SD(reg_array_23_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_24_) );
  senrq1 reg_array_reg_7__23_ ( .D(N775), .SD(reg_array_22_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_23_) );
  senrq1 reg_array_reg_7__22_ ( .D(N773), .SD(reg_array_21_), .ENN(n462), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_22_) );
  senrq1 reg_array_reg_7__21_ ( .D(N771), .SD(reg_array_20_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_21_) );
  senrq1 reg_array_reg_7__20_ ( .D(N769), .SD(reg_array_19_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_20_) );
  senrq1 reg_array_reg_7__19_ ( .D(N767), .SD(reg_array_18_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_19_) );
  senrq1 reg_array_reg_7__18_ ( .D(N765), .SD(reg_array_17_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_18_) );
  senrq1 reg_array_reg_7__17_ ( .D(N763), .SD(reg_array_16_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_17_) );
  senrq1 reg_array_reg_7__16_ ( .D(N761), .SD(reg_array_15_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_16_) );
  senrq1 reg_array_reg_7__15_ ( .D(N759), .SD(reg_array_14_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_15_) );
  senrq1 reg_array_reg_7__14_ ( .D(N757), .SD(reg_array_13_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_14_) );
  senrq1 reg_array_reg_7__13_ ( .D(N755), .SD(reg_array_12_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_13_) );
  senrq1 reg_array_reg_7__12_ ( .D(N753), .SD(reg_array_11_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_12_) );
  senrq1 reg_array_reg_7__11_ ( .D(N751), .SD(reg_array_10_), .ENN(n461), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_11_) );
  senrq1 reg_array_reg_7__10_ ( .D(N749), .SD(reg_array_9_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_10_) );
  senrq1 reg_array_reg_7__9_ ( .D(N747), .SD(reg_array_8_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_9_) );
  senrq1 reg_array_reg_7__8_ ( .D(N745), .SD(reg_array_7_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_8_) );
  senrq1 reg_array_reg_7__7_ ( .D(N743), .SD(reg_array_6_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_7_) );
  senrq1 reg_array_reg_7__6_ ( .D(N741), .SD(reg_array_5_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_6_) );
  senrq1 reg_array_reg_7__5_ ( .D(N739), .SD(reg_array_4_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_5_) );
  senrq1 reg_array_reg_7__4_ ( .D(N737), .SD(reg_array_3_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_4_) );
  senrq1 reg_array_reg_7__3_ ( .D(N735), .SD(reg_array_2_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_3_) );
  senrq1 reg_array_reg_7__2_ ( .D(N733), .SD(reg_array_1_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_2_) );
  senrq1 reg_array_reg_7__1_ ( .D(N731), .SD(reg_array_0_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_1_) );
  senrq1 reg_array_reg_7__0_ ( .D(N729), .SD(reg_array_63_), .ENN(n460), .SC(
        test_se), .CP(fifo_clk_push), .Q(reg_array_0_) );
  sdnrq1 data_out_reg_31_ ( .D(test_so1), .SD(data_out_fifo[30]), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_fifo[31]) );
  sdnrq1 data_out_reg_30_ ( .D(data_out_sync_30_), .SD(data_out_fifo[29]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[30]) );
  sdnrq1 data_out_reg_29_ ( .D(data_out_sync_29_), .SD(data_out_fifo[28]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[29]) );
  sdnrq1 data_out_reg_28_ ( .D(data_out_sync_28_), .SD(data_out_fifo[27]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[28]) );
  sdnrq1 data_out_reg_27_ ( .D(data_out_sync_27_), .SD(data_out_fifo[26]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[27]) );
  sdnrq1 data_out_reg_26_ ( .D(data_out_sync_26_), .SD(data_out_fifo[25]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[26]) );
  sdnrq1 data_out_reg_25_ ( .D(data_out_sync_25_), .SD(data_out_fifo[24]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[25]) );
  sdnrq1 data_out_reg_24_ ( .D(data_out_sync_24_), .SD(data_out_fifo[23]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[24]) );
  sdnrq1 data_out_reg_15_ ( .D(data_out_sync_15_), .SD(data_out_fifo[14]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[15]) );
  sdnrq1 data_out_reg_14_ ( .D(data_out_sync_14_), .SD(data_out_fifo[13]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[14]) );
  sdnrq1 data_out_reg_13_ ( .D(data_out_sync_13_), .SD(data_out_fifo[12]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[13]) );
  sdnrq1 data_out_reg_12_ ( .D(data_out_sync_12_), .SD(data_out_fifo[11]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[12]) );
  sdnrq1 data_out_reg_11_ ( .D(data_out_sync_11_), .SD(data_out_fifo[10]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[11]) );
  sdnrq1 data_out_reg_10_ ( .D(data_out_sync_10_), .SD(test_si1), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_fifo[10]) );
  sdnrq1 data_out_reg_9_ ( .D(data_out_sync_9_), .SD(data_out_fifo[8]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[9]) );
  sdnrq1 data_out_reg_8_ ( .D(data_out_sync_8_), .SD(data_out_fifo[7]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[8]) );
  sdnrq1 data_out_reg_23_ ( .D(data_out_sync_23_), .SD(data_out_fifo[22]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[23]) );
  sdnrq1 data_out_reg_22_ ( .D(data_out_sync_22_), .SD(data_out_fifo[21]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[22]) );
  sdnrq1 data_out_reg_21_ ( .D(data_out_sync_21_), .SD(data_out_fifo[20]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[21]) );
  sdnrq1 data_out_reg_20_ ( .D(data_out_sync_20_), .SD(data_out_fifo[19]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[20]) );
  sdnrq1 data_out_reg_19_ ( .D(data_out_sync_19_), .SD(data_out_fifo[18]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[19]) );
  sdnrq1 data_out_reg_18_ ( .D(data_out_sync_18_), .SD(data_out_fifo[17]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[18]) );
  sdnrq1 data_out_reg_17_ ( .D(data_out_sync_17_), .SD(data_out_fifo[16]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[17]) );
  sdnrq1 data_out_reg_16_ ( .D(data_out_sync_16_), .SD(data_out_fifo[15]), 
        .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[16]) );
  sdnrq1 data_out_reg_6_ ( .D(data_out_sync_6_), .SD(data_out_fifo[5]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[6]) );
  sdnrq1 data_out_reg_5_ ( .D(data_out_sync_5_), .SD(data_out_fifo[4]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[5]) );
  sdnrq1 data_out_reg_4_ ( .D(data_out_sync_4_), .SD(data_out_fifo[3]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[4]) );
  sdnrq1 data_out_reg_3_ ( .D(data_out_sync_3_), .SD(data_out_fifo[2]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[3]) );
  sdnrq1 data_out_reg_2_ ( .D(data_out_sync_2_), .SD(data_out_fifo[1]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[2]) );
  sdnrq1 data_out_reg_1_ ( .D(data_out_sync_1_), .SD(data_out_fifo[0]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[1]) );
  sdnrq1 data_out_reg_0_ ( .D(data_out_sync_0_), .SD(n465), .SC(test_se), .CP(
        fifo_clk_pop), .Q(data_out_fifo[0]) );
  sdnrq1 data_out_reg_7_ ( .D(data_out_sync_7_), .SD(data_out_fifo[6]), .SC(
        test_se), .CP(fifo_clk_pop), .Q(data_out_fifo[7]) );
  sdnrq1 data_out_sync_reg_31_ ( .D(N807), .SD(data_out_sync_30_), .SC(test_se), .CP(fifo_clk_pop), .Q(test_so1) );
  sdnrq1 data_out_sync_reg_30_ ( .D(N808), .SD(data_out_sync_29_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_30_) );
  sdnrq1 data_out_sync_reg_29_ ( .D(N809), .SD(data_out_sync_28_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_29_) );
  sdnrq1 data_out_sync_reg_28_ ( .D(N810), .SD(data_out_sync_27_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_28_) );
  sdnrq1 data_out_sync_reg_27_ ( .D(N811), .SD(data_out_sync_26_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_27_) );
  sdnrq1 data_out_sync_reg_26_ ( .D(N812), .SD(data_out_sync_25_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_26_) );
  sdnrq1 data_out_sync_reg_25_ ( .D(N813), .SD(data_out_sync_24_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_25_) );
  sdnrq1 data_out_sync_reg_24_ ( .D(N814), .SD(data_out_sync_23_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_24_) );
  sdnrq1 data_out_sync_reg_23_ ( .D(N815), .SD(data_out_sync_22_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_23_) );
  sdnrq1 data_out_sync_reg_22_ ( .D(N816), .SD(data_out_sync_21_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_22_) );
  sdnrq1 data_out_sync_reg_21_ ( .D(N817), .SD(data_out_sync_20_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_21_) );
  sdnrq1 data_out_sync_reg_20_ ( .D(N818), .SD(data_out_sync_19_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_20_) );
  sdnrq1 data_out_sync_reg_19_ ( .D(N819), .SD(data_out_sync_18_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_19_) );
  sdnrq1 data_out_sync_reg_18_ ( .D(N820), .SD(data_out_sync_17_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_18_) );
  sdnrq1 data_out_sync_reg_17_ ( .D(N821), .SD(data_out_sync_16_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_17_) );
  sdnrq1 data_out_sync_reg_16_ ( .D(N822), .SD(data_out_sync_15_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_16_) );
  sdnrq1 data_out_sync_reg_15_ ( .D(N823), .SD(data_out_sync_14_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_15_) );
  sdnrq1 data_out_sync_reg_14_ ( .D(N824), .SD(data_out_sync_13_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_14_) );
  sdnrq1 data_out_sync_reg_13_ ( .D(N825), .SD(data_out_sync_12_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_13_) );
  sdnrq1 data_out_sync_reg_12_ ( .D(N826), .SD(data_out_sync_11_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_12_) );
  sdnrq1 data_out_sync_reg_11_ ( .D(N827), .SD(data_out_sync_10_), .SC(test_se), .CP(fifo_clk_pop), .Q(data_out_sync_11_) );
  sdnrq1 data_out_sync_reg_10_ ( .D(N828), .SD(data_out_sync_9_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_10_) );
  sdnrq1 data_out_sync_reg_9_ ( .D(N829), .SD(data_out_sync_8_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_9_) );
  sdnrq1 data_out_sync_reg_8_ ( .D(N830), .SD(data_out_sync_7_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_8_) );
  sdnrq1 data_out_sync_reg_7_ ( .D(N831), .SD(data_out_sync_6_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_7_) );
  sdnrq1 data_out_sync_reg_6_ ( .D(N832), .SD(data_out_sync_5_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_6_) );
  sdnrq1 data_out_sync_reg_5_ ( .D(N833), .SD(data_out_sync_4_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_5_) );
  sdnrq1 data_out_sync_reg_4_ ( .D(N834), .SD(data_out_sync_3_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_4_) );
  sdnrq1 data_out_sync_reg_3_ ( .D(N835), .SD(data_out_sync_2_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_3_) );
  sdnrq1 data_out_sync_reg_2_ ( .D(N836), .SD(data_out_sync_1_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_2_) );
  sdnrq1 data_out_sync_reg_1_ ( .D(N837), .SD(data_out_sync_0_), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_1_) );
  sdnrq1 data_out_sync_reg_0_ ( .D(N838), .SD(data_out_fifo[31]), .SC(test_se), 
        .CP(fifo_clk_pop), .Q(data_out_sync_0_) );
  inv0d1 U98 ( .I(we_n), .ZN(n406) );
  bufbd1 U131 ( .I(n337), .Z(n422) );
  bufbd1 U164 ( .I(n337), .Z(n421) );
  bufbd1 U197 ( .I(n97), .Z(n460) );
  bufbd1 U230 ( .I(n97), .Z(n461) );
  bufbd1 U263 ( .I(n130), .Z(n457) );
  bufbd1 U296 ( .I(n130), .Z(n458) );
  bufbd1 U329 ( .I(n163), .Z(n454) );
  bufbd1 U331 ( .I(n163), .Z(n455) );
  bufbd1 U332 ( .I(n1), .Z(n451) );
  bufbd1 U333 ( .I(n1), .Z(n452) );
  bufbd1 U334 ( .I(n196), .Z(n448) );
  bufbd1 U335 ( .I(n196), .Z(n449) );
  bufbd1 U336 ( .I(n229), .Z(n445) );
  bufbd1 U337 ( .I(n229), .Z(n446) );
  bufbd1 U338 ( .I(n262), .Z(n442) );
  bufbd1 U339 ( .I(n262), .Z(n443) );
  bufbd1 U340 ( .I(n295), .Z(n439) );
  bufbd1 U341 ( .I(n295), .Z(n440) );
  bufbd1 U342 ( .I(n337), .Z(n423) );
  bufbd1 U343 ( .I(n97), .Z(n462) );
  bufbd1 U344 ( .I(n130), .Z(n459) );
  bufbd1 U345 ( .I(n163), .Z(n456) );
  bufbd1 U346 ( .I(n1), .Z(n453) );
  bufbd1 U347 ( .I(n196), .Z(n450) );
  bufbd1 U348 ( .I(n229), .Z(n447) );
  bufbd1 U349 ( .I(n262), .Z(n444) );
  bufbd1 U350 ( .I(n295), .Z(n441) );
  bufbd1 U351 ( .I(n339), .Z(n416) );
  bufbd1 U352 ( .I(n336), .Z(n425) );
  bufbd1 U353 ( .I(n338), .Z(n419) );
  bufbd1 U354 ( .I(n339), .Z(n404) );
  bufbd1 U355 ( .I(n336), .Z(n424) );
  bufbd1 U356 ( .I(n338), .Z(n418) );
  bufbd1 U357 ( .I(n339), .Z(n417) );
  bufbd1 U358 ( .I(n336), .Z(n426) );
  bufbd1 U359 ( .I(n338), .Z(n420) );
  bufbd1 U360 ( .I(n333), .Z(n434) );
  bufbd1 U361 ( .I(n335), .Z(n428) );
  bufbd1 U362 ( .I(n334), .Z(n431) );
  bufbd1 U367 ( .I(n332), .Z(n437) );
  bufbd1 U368 ( .I(n333), .Z(n433) );
  bufbd1 U369 ( .I(n335), .Z(n427) );
  bufbd1 U370 ( .I(n334), .Z(n430) );
  bufbd1 U371 ( .I(n332), .Z(n436) );
  bufbd1 U372 ( .I(n333), .Z(n435) );
  bufbd1 U373 ( .I(n335), .Z(n429) );
  bufbd1 U374 ( .I(n334), .Z(n432) );
  bufbd1 U375 ( .I(n332), .Z(n438) );
  an02d1 U376 ( .A1(fifo_rst_n), .A2(n412), .Z(n1) );
  inv0d1 U377 ( .I(rd_addr[1]), .ZN(n403) );
  inv0d1 U378 ( .I(wr_addr[1]), .ZN(n407) );
  inv0d1 U411 ( .I(wr_addr[2]), .ZN(n408) );
  an02d1 U412 ( .A1(fifo_rst_n), .A2(n415), .Z(n97) );
  an02d1 U481 ( .A1(fifo_rst_n), .A2(n414), .Z(n130) );
  an02d1 U489 ( .A1(fifo_rst_n), .A2(n413), .Z(n163) );
  an02d1 U490 ( .A1(fifo_rst_n), .A2(n411), .Z(n196) );
  an02d1 U491 ( .A1(fifo_rst_n), .A2(n409), .Z(n229) );
  inv0d1 U492 ( .I(wr_addr[0]), .ZN(n410) );
  an02d1 U493 ( .A1(fifo_rst_n), .A2(n405), .Z(n262) );
  an02d1 U494 ( .A1(n328), .A2(fifo_rst_n), .Z(n295) );
  or04d1 U495 ( .A1(wr_addr[2]), .A2(wr_addr[1]), .A3(wr_addr[0]), .A4(we_n), 
        .Z(n328) );
  nd02d1 U496 ( .A1(n330), .A2(n331), .ZN(N838) );
  nd02d1 U497 ( .A1(n340), .A2(n341), .ZN(N837) );
  nd02d1 U498 ( .A1(n342), .A2(n343), .ZN(N836) );
  nd02d1 U499 ( .A1(n344), .A2(n345), .ZN(N835) );
  nd02d1 U500 ( .A1(n346), .A2(n347), .ZN(N834) );
  nd02d1 U501 ( .A1(n348), .A2(n349), .ZN(N833) );
  nd02d1 U502 ( .A1(n350), .A2(n351), .ZN(N832) );
  nd02d1 U503 ( .A1(n352), .A2(n353), .ZN(N831) );
  nd02d1 U504 ( .A1(n354), .A2(n355), .ZN(N830) );
  nd02d1 U505 ( .A1(n356), .A2(n357), .ZN(N829) );
  nd02d1 U506 ( .A1(n358), .A2(n359), .ZN(N828) );
  nd02d1 U507 ( .A1(n360), .A2(n361), .ZN(N827) );
  nd02d1 U508 ( .A1(n362), .A2(n363), .ZN(N826) );
  nd02d1 U509 ( .A1(n364), .A2(n365), .ZN(N825) );
  nd02d1 U510 ( .A1(n366), .A2(n367), .ZN(N824) );
  nd02d1 U511 ( .A1(n368), .A2(n369), .ZN(N823) );
  nd02d1 U512 ( .A1(n370), .A2(n371), .ZN(N822) );
  nd02d1 U513 ( .A1(n372), .A2(n373), .ZN(N821) );
  nd02d1 U514 ( .A1(n374), .A2(n375), .ZN(N820) );
  nd02d1 U515 ( .A1(n376), .A2(n377), .ZN(N819) );
  nd02d1 U516 ( .A1(n378), .A2(n379), .ZN(N818) );
  nd02d1 U517 ( .A1(n380), .A2(n381), .ZN(N817) );
  nd02d1 U518 ( .A1(n382), .A2(n383), .ZN(N816) );
  nd02d1 U519 ( .A1(n384), .A2(n385), .ZN(N815) );
  nd02d1 U520 ( .A1(n386), .A2(n387), .ZN(N814) );
  nd02d1 U521 ( .A1(n388), .A2(n389), .ZN(N813) );
  nd02d1 U522 ( .A1(n390), .A2(n391), .ZN(N812) );
  nd02d1 U523 ( .A1(n392), .A2(n393), .ZN(N811) );
  nd02d1 U524 ( .A1(n394), .A2(n395), .ZN(N810) );
  nd02d1 U525 ( .A1(n396), .A2(n397), .ZN(N809) );
  nd02d1 U526 ( .A1(n398), .A2(n399), .ZN(N808) );
  nd02d1 U527 ( .A1(n400), .A2(n401), .ZN(N807) );
  inv0d1 U528 ( .I(rd_addr[0]), .ZN(n402) );
endmodule


module SDRAM_IF ( sdram_clk, sdram_rst_n, risc_OUT_VALID, risc_STACK_FULL, 
        risc_EndOfInstrn, risc_PSW, risc_Rd_Instr, sd_A, sd_CK, sd_CKn, sd_LD, 
        sd_RW, sd_BWS, sd_DQ_in, sd_DQ_out, sd_DQ_en, sd_wfifo_pop, 
        sd_wfifo_empty, sd_rfifo_push, sd_rfifo_full, sd_rfifo_DQ_out, 
        sd_wfifo_DQ_in, test_se, test_si1, test_si2, test_si3, test_so2, 
        test_so1 );
  input [10:0] risc_PSW;
  output [9:0] sd_A;
  output [1:0] sd_BWS;
  input [15:0] sd_DQ_in;
  output [15:0] sd_DQ_out;
  output [15:0] sd_DQ_en;
  output [31:0] sd_rfifo_DQ_out;
  input [31:0] sd_wfifo_DQ_in;
  input sdram_clk, sdram_rst_n, risc_OUT_VALID, risc_STACK_FULL,
         risc_EndOfInstrn, risc_Rd_Instr, sd_wfifo_empty, sd_rfifo_full,
         test_se, test_si1, test_si2, test_si3;
  output sd_CK, sd_CKn, sd_LD, sd_RW, sd_wfifo_pop, sd_rfifo_push, test_so2,
         test_so1;
  wire   n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, N7, sync_control_bus_13_,
         sync_control_bus_12_, sync_control_bus_11_, sync_control_bus_10_,
         sync_control_bus_9_, sync_control_bus_8_, sync_control_bus_7_,
         sync_control_bus_6_, sync_control_bus_5_, sync_control_bus_4_,
         sync_control_bus_3_, sync_control_bus_2_, sync_control_bus_1_,
         sync_control_bus_0_, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N390, N630, N870, N990, mega_shift_1_79_, mega_shift_1_78_,
         mega_shift_1_77_, mega_shift_1_76_, mega_shift_1_75_,
         mega_shift_1_74_, mega_shift_1_73_, mega_shift_1_72_,
         mega_shift_1_71_, mega_shift_1_70_, mega_shift_1_69_,
         mega_shift_1_68_, mega_shift_1_67_, mega_shift_1_66_,
         mega_shift_1_65_, mega_shift_1_64_, mega_shift_1_63_,
         mega_shift_1_62_, mega_shift_1_61_, mega_shift_1_60_,
         mega_shift_1_59_, mega_shift_1_58_, mega_shift_1_57_,
         mega_shift_1_56_, mega_shift_1_55_, mega_shift_1_54_,
         mega_shift_1_53_, mega_shift_1_52_, mega_shift_1_51_,
         mega_shift_1_50_, mega_shift_1_49_, mega_shift_1_48_,
         mega_shift_1_47_, mega_shift_1_46_, mega_shift_1_45_,
         mega_shift_1_44_, mega_shift_1_43_, mega_shift_1_42_,
         mega_shift_1_41_, mega_shift_1_40_, mega_shift_1_39_,
         mega_shift_1_38_, mega_shift_1_37_, mega_shift_1_36_,
         mega_shift_1_35_, mega_shift_1_34_, mega_shift_1_33_,
         mega_shift_1_32_, mega_shift_1_31_, mega_shift_1_30_,
         mega_shift_1_29_, mega_shift_1_28_, mega_shift_1_27_,
         mega_shift_1_26_, mega_shift_1_25_, mega_shift_1_24_,
         mega_shift_1_23_, mega_shift_1_22_, mega_shift_1_21_,
         mega_shift_1_20_, mega_shift_1_19_, mega_shift_1_18_,
         mega_shift_1_17_, mega_shift_1_16_, mega_shift_1_14_,
         mega_shift_1_13_, mega_shift_1_12_, mega_shift_1_11_,
         mega_shift_1_10_, mega_shift_1_9_, mega_shift_1_8_, mega_shift_1_7_,
         mega_shift_1_6_, mega_shift_1_5_, mega_shift_1_4_, mega_shift_1_3_,
         mega_shift_1_2_, mega_shift_1_1_, mega_shift_1_0_, N1350, N1590,
         N1830, N2070, n297, n308, n315, n318, n321, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n364, n365, n366, n367, n368, n369, n370, n371, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, add_167_carry_3_, add_167_carry_4_, add_167_carry_5_,
         add_167_carry_6_, add_167_carry_7_, add_167_carry_8_,
         add_167_carry_9_, add_167_carry_10_, add_167_carry_11_,
         add_167_carry_12_, add_167_carry_13_, add_167_carry_14_,
         add_167_carry_15_, add_165_carry_3_, add_165_carry_4_,
         add_165_carry_5_, add_165_carry_6_, add_165_carry_7_,
         add_165_carry_8_, add_165_carry_9_, add_165_carry_10_,
         add_165_carry_11_, add_165_carry_12_, add_165_carry_13_,
         add_165_carry_14_, add_165_carry_15_, add_163_carry_3_,
         add_163_carry_4_, add_163_carry_5_, add_163_carry_6_,
         add_163_carry_7_, add_163_carry_8_, add_163_carry_9_,
         add_163_carry_10_, add_163_carry_11_, add_163_carry_12_,
         add_163_carry_13_, add_163_carry_14_, add_163_carry_15_,
         add_161_carry_3_, add_161_carry_4_, add_161_carry_5_,
         add_161_carry_6_, add_161_carry_7_, add_161_carry_8_,
         add_161_carry_9_, add_161_carry_10_, add_161_carry_11_,
         add_161_carry_12_, add_161_carry_13_, add_161_carry_14_,
         add_161_carry_15_, add_159_carry_3_, add_159_carry_4_,
         add_159_carry_5_, add_159_carry_6_, add_159_carry_7_,
         add_159_carry_8_, add_159_carry_9_, add_159_carry_10_,
         add_159_carry_11_, add_159_carry_12_, add_159_carry_13_,
         add_159_carry_14_, add_159_carry_15_, add_157_carry_4_,
         add_157_carry_5_, add_157_carry_6_, add_157_carry_7_,
         add_157_carry_8_, add_157_carry_9_, add_157_carry_10_,
         add_157_carry_11_, add_157_carry_12_, add_157_carry_13_,
         add_157_carry_14_, add_157_carry_15_, add_155_carry_6_,
         add_155_carry_7_, add_155_carry_8_, add_155_carry_9_,
         add_155_carry_10_, add_155_carry_11_, add_155_carry_12_,
         add_155_carry_13_, add_155_carry_14_, add_155_carry_15_,
         add_153_carry_3_, add_153_carry_4_, add_153_carry_5_,
         add_153_carry_6_, add_153_carry_7_, add_153_carry_8_,
         add_153_carry_9_, add_153_carry_10_, add_153_carry_11_,
         add_153_carry_12_, add_153_carry_13_, add_153_carry_14_,
         add_153_carry_15_, n17, n363, n372, n383, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518;
  wire   [15:0] c_out_control;
  wire   [14:0] control_bus;
  wire   [79:0] mega_shift_0;
  wire   [15:0] DQ_out_0;
  wire   [15:0] DQ_out_1;

  mx02d4 sd_mux_dq_out_15 ( .I0(DQ_out_0[15]), .I1(DQ_out_1[15]), .S(sdram_clk), .Z(sd_DQ_out[15]) );
  mx02d4 sd_mux_dq_out_14 ( .I0(DQ_out_0[14]), .I1(DQ_out_1[14]), .S(sdram_clk), .Z(sd_DQ_out[14]) );
  mx02d4 sd_mux_dq_out_13 ( .I0(DQ_out_0[13]), .I1(DQ_out_1[13]), .S(sdram_clk), .Z(sd_DQ_out[13]) );
  mx02d4 sd_mux_dq_out_12 ( .I0(DQ_out_0[12]), .I1(DQ_out_1[12]), .S(sdram_clk), .Z(sd_DQ_out[12]) );
  mx02d4 sd_mux_dq_out_11 ( .I0(DQ_out_0[11]), .I1(DQ_out_1[11]), .S(sdram_clk), .Z(sd_DQ_out[11]) );
  mx02d4 sd_mux_dq_out_10 ( .I0(DQ_out_0[10]), .I1(DQ_out_1[10]), .S(sdram_clk), .Z(sd_DQ_out[10]) );
  mx02d4 sd_mux_dq_out_9 ( .I0(DQ_out_0[9]), .I1(DQ_out_1[9]), .S(sdram_clk), 
        .Z(sd_DQ_out[9]) );
  mx02d4 sd_mux_dq_out_8 ( .I0(DQ_out_0[8]), .I1(DQ_out_1[8]), .S(sdram_clk), 
        .Z(sd_DQ_out[8]) );
  mx02d4 sd_mux_dq_out_7 ( .I0(DQ_out_0[7]), .I1(DQ_out_1[7]), .S(sdram_clk), 
        .Z(sd_DQ_out[7]) );
  mx02d4 sd_mux_dq_out_6 ( .I0(DQ_out_0[6]), .I1(DQ_out_1[6]), .S(sdram_clk), 
        .Z(sd_DQ_out[6]) );
  mx02d4 sd_mux_dq_out_5 ( .I0(DQ_out_0[5]), .I1(DQ_out_1[5]), .S(sdram_clk), 
        .Z(sd_DQ_out[5]) );
  mx02d4 sd_mux_dq_out_4 ( .I0(DQ_out_0[4]), .I1(DQ_out_1[4]), .S(sdram_clk), 
        .Z(sd_DQ_out[4]) );
  mx02d4 sd_mux_dq_out_3 ( .I0(DQ_out_0[3]), .I1(DQ_out_1[3]), .S(sdram_clk), 
        .Z(sd_DQ_out[3]) );
  mx02d4 sd_mux_dq_out_2 ( .I0(DQ_out_0[2]), .I1(DQ_out_1[2]), .S(sdram_clk), 
        .Z(sd_DQ_out[2]) );
  mx02d4 sd_mux_dq_out_1 ( .I0(DQ_out_0[1]), .I1(DQ_out_1[1]), .S(sdram_clk), 
        .Z(sd_DQ_out[1]) );
  mx02d4 sd_mux_dq_out_0 ( .I0(DQ_out_0[0]), .I1(DQ_out_1[0]), .S(sdram_clk), 
        .Z(sd_DQ_out[0]) );
  mx02d4 sd_mux_CK ( .I0(1'b0), .I1(1'b1), .S(sdram_clk), .Z(sd_CK) );
  mx02d4 sd_mux_CKn ( .I0(1'b1), .I1(1'b0), .S(sdram_clk), .Z(sd_CKn) );
  sdnrn1 control_bus_reg_13_ ( .D(sync_control_bus_13_), .SD(control_bus[12]), 
        .SC(test_se), .CP(sdram_clk), .QN(n321) );
  sdnrn1 control_bus_reg_12_ ( .D(sync_control_bus_12_), .SD(control_bus[11]), 
        .SC(test_se), .CP(sdram_clk), .QN(n318) );
  sdnrn1 control_bus_reg_11_ ( .D(sync_control_bus_11_), .SD(n479), .SC(
        test_se), .CP(sdram_clk), .QN(n315) );
  sdnrn1 control_bus_reg_8_ ( .D(sync_control_bus_8_), .SD(n475), .SC(test_se), 
        .CP(sdram_clk), .QN(n308) );
  sdnrn1 control_bus_reg_3_ ( .D(sync_control_bus_3_), .SD(N43), .SC(test_se), 
        .CP(sdram_clk), .QN(n297) );
  sdnfb1 DQ_in_1_reg_15_ ( .D(sd_DQ_in[15]), .SD(n504), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[31]), .QN(n503) );
  sdnfb1 DQ_in_1_reg_14_ ( .D(sd_DQ_in[14]), .SD(n505), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[30]), .QN(n504) );
  sdnfb1 DQ_in_1_reg_13_ ( .D(sd_DQ_in[13]), .SD(n506), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[29]), .QN(n505) );
  sdnfb1 DQ_in_1_reg_12_ ( .D(sd_DQ_in[12]), .SD(n507), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[28]), .QN(n506) );
  sdnfb1 DQ_in_1_reg_11_ ( .D(sd_DQ_in[11]), .SD(n508), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[27]), .QN(n507) );
  sdnfb1 DQ_in_1_reg_10_ ( .D(sd_DQ_in[10]), .SD(n509), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[26]), .QN(n508) );
  sdnfb1 DQ_in_1_reg_9_ ( .D(sd_DQ_in[9]), .SD(n510), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[25]), .QN(n509) );
  sdnfb1 DQ_in_1_reg_8_ ( .D(sd_DQ_in[8]), .SD(n511), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[24]), .QN(n510) );
  sdnfb1 DQ_in_1_reg_7_ ( .D(sd_DQ_in[7]), .SD(n512), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[23]), .QN(n511) );
  sdnfb1 DQ_in_1_reg_6_ ( .D(sd_DQ_in[6]), .SD(n513), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[22]), .QN(n512) );
  sdnfb1 DQ_in_1_reg_5_ ( .D(sd_DQ_in[5]), .SD(n514), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[21]), .QN(n513) );
  sdnfb1 DQ_in_1_reg_4_ ( .D(sd_DQ_in[4]), .SD(n515), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[20]), .QN(n514) );
  sdnfb1 DQ_in_1_reg_3_ ( .D(sd_DQ_in[3]), .SD(n516), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[19]), .QN(n515) );
  sdnfb1 DQ_in_1_reg_2_ ( .D(sd_DQ_in[2]), .SD(n517), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[18]), .QN(n516) );
  sdnfb1 DQ_in_1_reg_1_ ( .D(sd_DQ_in[1]), .SD(n518), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[17]), .QN(n517) );
  sdnfb1 DQ_in_1_reg_0_ ( .D(sd_DQ_in[0]), .SD(test_si2), .SC(test_se), .CPN(
        sdram_clk), .Q(sd_rfifo_DQ_out[16]), .QN(n518) );
  an04d1 U323 ( .A1(n371), .A2(n315), .A3(n373), .A4(n374), .Z(n370) );
  an03d1 U330 ( .A1(n383), .A2(n381), .A3(n472), .Z(n389) );
  an03d1 U331 ( .A1(control_bus[12]), .A2(n376), .A3(n390), .Z(n381) );
  an03d1 U332 ( .A1(control_bus[4]), .A2(n481), .A3(n483), .Z(n376) );
  an03d1 U333 ( .A1(N42), .A2(n391), .A3(control_bus[9]), .Z(n386) );
  an03d1 U334 ( .A1(n477), .A2(control_bus[3]), .A3(n392), .Z(n373) );
  an04d1 U339 ( .A1(n469), .A2(control_bus[14]), .A3(n369), .A4(n297), .Z(n375) );
  aoi2222d1 U382 ( .A1(N143), .A2(n327), .B1(N127), .B2(n328), .C1(N111), .C2(
        n329), .D1(N95), .D2(n330), .ZN(n326) );
  aoi2222d1 U383 ( .A1(N79), .A2(n331), .B1(N63), .B2(n332), .C1(N47), .C2(
        n333), .D1(N31), .D2(n334), .ZN(n325) );
  aoi2222d1 U384 ( .A1(N142), .A2(n327), .B1(N126), .B2(n328), .C1(N110), .C2(
        n329), .D1(N94), .D2(n330), .ZN(n336) );
  aoi2222d1 U385 ( .A1(N78), .A2(n331), .B1(N62), .B2(n332), .C1(N46), .C2(
        n333), .D1(N30), .D2(n334), .ZN(n335) );
  aoi2222d1 U386 ( .A1(N141), .A2(n327), .B1(N125), .B2(n328), .C1(N109), .C2(
        n329), .D1(N93), .D2(n330), .ZN(n338) );
  aoi2222d1 U387 ( .A1(N77), .A2(n331), .B1(N61), .B2(n332), .C1(N45), .C2(
        n333), .D1(N29), .D2(n334), .ZN(n337) );
  aoi2222d1 U388 ( .A1(N140), .A2(n327), .B1(N124), .B2(n328), .C1(N108), .C2(
        n329), .D1(N92), .D2(n330), .ZN(n340) );
  aoi2222d1 U389 ( .A1(N76), .A2(n331), .B1(N60), .B2(n332), .C1(N44), .C2(
        n333), .D1(N28), .D2(n334), .ZN(n339) );
  aoi2222d1 U390 ( .A1(N139), .A2(n327), .B1(N123), .B2(n328), .C1(N107), .C2(
        n329), .D1(N91), .D2(n330), .ZN(n342) );
  aoi2222d1 U391 ( .A1(N75), .A2(n331), .B1(N59), .B2(n332), .C1(N43), .C2(
        n333), .D1(N27), .D2(n334), .ZN(n341) );
  aoi2222d1 U392 ( .A1(N138), .A2(n327), .B1(N122), .B2(n328), .C1(N106), .C2(
        n329), .D1(N90), .D2(n330), .ZN(n344) );
  aoi2222d1 U393 ( .A1(N74), .A2(n331), .B1(N58), .B2(n332), .C1(N42), .C2(
        n333), .D1(N26), .D2(n334), .ZN(n343) );
  aoi2222d1 U394 ( .A1(N137), .A2(n327), .B1(N121), .B2(n328), .C1(N105), .C2(
        n329), .D1(N89), .D2(n330), .ZN(n346) );
  aoi2222d1 U395 ( .A1(N73), .A2(n331), .B1(N57), .B2(n332), .C1(n363), .C2(
        n333), .D1(N25), .D2(n334), .ZN(n345) );
  aoi2222d1 U396 ( .A1(N136), .A2(n327), .B1(N120), .B2(n328), .C1(N104), .C2(
        n329), .D1(N88), .D2(n330), .ZN(n348) );
  aoi2222d1 U397 ( .A1(N72), .A2(n331), .B1(N56), .B2(n332), .C1(n482), .C2(
        n333), .D1(N24), .D2(n334), .ZN(n347) );
  aoi2222d1 U398 ( .A1(N23), .A2(n327), .B1(N23), .B2(n328), .C1(N23), .C2(
        n329), .D1(N23), .D2(n330), .ZN(n350) );
  aoi2222d1 U399 ( .A1(N23), .A2(n331), .B1(n483), .B2(n332), .C1(n483), .C2(
        n333), .D1(N23), .D2(n334), .ZN(n349) );
  aoi2222d1 U400 ( .A1(N149), .A2(n327), .B1(N133), .B2(n328), .C1(N117), .C2(
        n329), .D1(N101), .D2(n330), .ZN(n352) );
  aoi2222d1 U401 ( .A1(N85), .A2(n331), .B1(N69), .B2(n332), .C1(N53), .C2(
        n333), .D1(N37), .D2(n334), .ZN(n351) );
  aoi2222d1 U402 ( .A1(N148), .A2(n327), .B1(N132), .B2(n328), .C1(N116), .C2(
        n329), .D1(N100), .D2(n330), .ZN(n354) );
  aoi2222d1 U403 ( .A1(N84), .A2(n331), .B1(N68), .B2(n332), .C1(N52), .C2(
        n333), .D1(N36), .D2(n334), .ZN(n353) );
  aoi2222d1 U404 ( .A1(N147), .A2(n327), .B1(N131), .B2(n328), .C1(N115), .C2(
        n329), .D1(N99), .D2(n330), .ZN(n356) );
  aoi2222d1 U405 ( .A1(N83), .A2(n331), .B1(N67), .B2(n332), .C1(N51), .C2(
        n333), .D1(N35), .D2(n334), .ZN(n355) );
  aoi2222d1 U406 ( .A1(N146), .A2(n327), .B1(N130), .B2(n328), .C1(N114), .C2(
        n329), .D1(N98), .D2(n330), .ZN(n358) );
  aoi2222d1 U407 ( .A1(N82), .A2(n331), .B1(N66), .B2(n332), .C1(N50), .C2(
        n333), .D1(N34), .D2(n334), .ZN(n357) );
  aoi2222d1 U408 ( .A1(N145), .A2(n327), .B1(N129), .B2(n328), .C1(N113), .C2(
        n329), .D1(N97), .D2(n330), .ZN(n360) );
  aoi2222d1 U409 ( .A1(N81), .A2(n331), .B1(N65), .B2(n332), .C1(N49), .C2(
        n333), .D1(N33), .D2(n334), .ZN(n359) );
  aoi2222d1 U410 ( .A1(N144), .A2(n327), .B1(N128), .B2(n328), .C1(N112), .C2(
        n329), .D1(N96), .D2(n330), .ZN(n362) );
  aoi2222d1 U411 ( .A1(N80), .A2(n331), .B1(N64), .B2(n332), .C1(N48), .C2(
        n333), .D1(N32), .D2(n334), .ZN(n361) );
  nr04d0 U413 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(n368) );
  nd04d0 U414 ( .A1(n480), .A2(n369), .A3(n372), .A4(n370), .ZN(n367) );
  nd04d0 U415 ( .A1(n375), .A2(n376), .A3(n377), .A4(n378), .ZN(n365) );
  nr03d0 U416 ( .A1(n315), .A2(n379), .A3(n380), .ZN(n378) );
  nd04d0 U417 ( .A1(n381), .A2(control_bus[14]), .A3(n377), .A4(n382), .ZN(
        n366) );
  nr04d0 U418 ( .A1(n476), .A2(n468), .A3(n297), .A4(n384), .ZN(n382) );
  nr04d0 U419 ( .A1(n371), .A2(n385), .A3(n372), .A4(n473), .ZN(n377) );
  nr03d0 U421 ( .A1(control_bus[11]), .A2(n482), .A3(control_bus[5]), .ZN(n390) );
  nr03d0 U422 ( .A1(n385), .A2(n469), .A3(control_bus[14]), .ZN(n392) );
  nr03d0 U423 ( .A1(n383), .A2(n481), .A3(n315), .ZN(n387) );
  nr04d0 U424 ( .A1(n379), .A2(control_bus[4]), .A3(n472), .A4(n483), .ZN(n374) );
  nd03d0 U425 ( .A1(control_bus[5]), .A2(n393), .A3(n482), .ZN(n379) );
  nr03d0 U426 ( .A1(N42), .A2(n476), .A3(control_bus[13]), .ZN(n388) );
  nr02d0 U427 ( .A1(n391), .A2(control_bus[9]), .ZN(n369) );
  xn02d1 U428 ( .A1(mega_shift_0[29]), .A2(mega_shift_0[28]), .ZN(n397) );
  xr02d1 U429 ( .A1(mega_shift_0[25]), .A2(mega_shift_0[24]), .Z(n398) );
  xn02d1 U430 ( .A1(n399), .A2(n400), .ZN(n394) );
  xr02d1 U431 ( .A1(mega_shift_0[19]), .A2(mega_shift_0[18]), .Z(n401) );
  xr02d1 U432 ( .A1(mega_shift_0[23]), .A2(mega_shift_0[22]), .Z(n402) );
  xn02d1 U433 ( .A1(mega_shift_0[45]), .A2(mega_shift_0[44]), .ZN(n406) );
  xr02d1 U434 ( .A1(mega_shift_0[41]), .A2(mega_shift_0[40]), .Z(n407) );
  xn02d1 U435 ( .A1(n408), .A2(n409), .ZN(n403) );
  xr02d1 U436 ( .A1(mega_shift_0[35]), .A2(mega_shift_0[34]), .Z(n410) );
  xr02d1 U437 ( .A1(mega_shift_0[39]), .A2(mega_shift_0[38]), .Z(n411) );
  xn02d1 U438 ( .A1(mega_shift_1_13_), .A2(mega_shift_1_12_), .ZN(n415) );
  xr02d1 U439 ( .A1(mega_shift_1_9_), .A2(mega_shift_1_8_), .Z(n416) );
  xn02d1 U440 ( .A1(n417), .A2(n418), .ZN(n412) );
  xr02d1 U441 ( .A1(mega_shift_1_3_), .A2(mega_shift_1_2_), .Z(n419) );
  xr02d1 U442 ( .A1(mega_shift_1_7_), .A2(mega_shift_1_6_), .Z(n420) );
  xn02d1 U443 ( .A1(mega_shift_0[61]), .A2(mega_shift_0[60]), .ZN(n424) );
  xr02d1 U444 ( .A1(mega_shift_0[57]), .A2(mega_shift_0[56]), .Z(n425) );
  xn02d1 U445 ( .A1(n426), .A2(n427), .ZN(n421) );
  xr02d1 U446 ( .A1(mega_shift_0[51]), .A2(mega_shift_0[50]), .Z(n428) );
  xr02d1 U447 ( .A1(mega_shift_0[55]), .A2(mega_shift_0[54]), .Z(n429) );
  xn02d1 U448 ( .A1(mega_shift_1_29_), .A2(mega_shift_1_28_), .ZN(n433) );
  xr02d1 U449 ( .A1(mega_shift_1_25_), .A2(mega_shift_1_24_), .Z(n434) );
  xn02d1 U450 ( .A1(n435), .A2(n436), .ZN(n430) );
  xr02d1 U451 ( .A1(mega_shift_1_19_), .A2(mega_shift_1_18_), .Z(n437) );
  xr02d1 U452 ( .A1(mega_shift_1_23_), .A2(mega_shift_1_22_), .Z(n438) );
  xn02d1 U453 ( .A1(mega_shift_1_45_), .A2(mega_shift_1_44_), .ZN(n442) );
  xr02d1 U454 ( .A1(mega_shift_1_41_), .A2(mega_shift_1_40_), .Z(n443) );
  xn02d1 U455 ( .A1(n444), .A2(n445), .ZN(n439) );
  xr02d1 U456 ( .A1(mega_shift_1_35_), .A2(mega_shift_1_34_), .Z(n446) );
  xr02d1 U457 ( .A1(mega_shift_1_39_), .A2(mega_shift_1_38_), .Z(n447) );
  xn02d1 U458 ( .A1(mega_shift_1_61_), .A2(mega_shift_1_60_), .ZN(n451) );
  xr02d1 U459 ( .A1(mega_shift_1_57_), .A2(mega_shift_1_56_), .Z(n452) );
  xn02d1 U460 ( .A1(n453), .A2(n454), .ZN(n448) );
  xr02d1 U461 ( .A1(mega_shift_1_51_), .A2(mega_shift_1_50_), .Z(n455) );
  xr02d1 U462 ( .A1(mega_shift_1_55_), .A2(mega_shift_1_54_), .Z(n456) );
  xn02d1 U463 ( .A1(mega_shift_0[13]), .A2(mega_shift_0[12]), .ZN(n460) );
  xr02d1 U464 ( .A1(mega_shift_0[9]), .A2(mega_shift_0[8]), .Z(n461) );
  xn02d1 U465 ( .A1(n462), .A2(n463), .ZN(n457) );
  xr02d1 U466 ( .A1(mega_shift_0[3]), .A2(mega_shift_0[2]), .Z(n464) );
  xr02d1 U467 ( .A1(mega_shift_0[7]), .A2(mega_shift_0[6]), .Z(n465) );
  sdnrq1 DQ_in_0_reg_15_ ( .D(sd_DQ_in[15]), .SD(sd_rfifo_DQ_out[14]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[15]) );
  sdnrq1 DQ_in_0_reg_14_ ( .D(sd_DQ_in[14]), .SD(sd_rfifo_DQ_out[13]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[14]) );
  sdnrq1 DQ_in_0_reg_13_ ( .D(sd_DQ_in[13]), .SD(sd_rfifo_DQ_out[12]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[13]) );
  sdnrq1 DQ_in_0_reg_12_ ( .D(sd_DQ_in[12]), .SD(sd_rfifo_DQ_out[11]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[12]) );
  sdnrq1 DQ_in_0_reg_11_ ( .D(sd_DQ_in[11]), .SD(sd_rfifo_DQ_out[10]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[11]) );
  sdnrq1 DQ_in_0_reg_10_ ( .D(sd_DQ_in[10]), .SD(sd_rfifo_DQ_out[9]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[10]) );
  sdnrq1 DQ_in_0_reg_9_ ( .D(sd_DQ_in[9]), .SD(sd_rfifo_DQ_out[8]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[9]) );
  sdnrq1 DQ_in_0_reg_8_ ( .D(sd_DQ_in[8]), .SD(sd_rfifo_DQ_out[7]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[8]) );
  sdnrq1 DQ_in_0_reg_7_ ( .D(sd_DQ_in[7]), .SD(sd_rfifo_DQ_out[6]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[7]) );
  sdnrq1 DQ_in_0_reg_6_ ( .D(sd_DQ_in[6]), .SD(sd_rfifo_DQ_out[5]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[6]) );
  sdnrq1 DQ_in_0_reg_5_ ( .D(sd_DQ_in[5]), .SD(sd_rfifo_DQ_out[4]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[5]) );
  sdnrq1 DQ_in_0_reg_4_ ( .D(sd_DQ_in[4]), .SD(sd_rfifo_DQ_out[3]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[4]) );
  sdnrq1 DQ_in_0_reg_3_ ( .D(sd_DQ_in[3]), .SD(sd_rfifo_DQ_out[2]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[3]) );
  sdnrq1 DQ_in_0_reg_2_ ( .D(sd_DQ_in[2]), .SD(sd_rfifo_DQ_out[1]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[2]) );
  sdnrq1 DQ_in_0_reg_1_ ( .D(sd_DQ_in[1]), .SD(sd_rfifo_DQ_out[0]), .SC(
        test_se), .CP(sdram_clk), .Q(sd_rfifo_DQ_out[1]) );
  sdnrq1 DQ_in_0_reg_0_ ( .D(sd_DQ_in[0]), .SD(test_si1), .SC(test_se), .CP(
        sdram_clk), .Q(sd_rfifo_DQ_out[0]) );
  sdcrq1 mega_shift_0_reg_4__15_ ( .D(sd_wfifo_DQ_in[15]), .SD(
        mega_shift_0[14]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_0[15]) );
  sdcrq1 mega_shift_0_reg_3__15_ ( .D(N990), .SD(mega_shift_0[30]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[31]) );
  sdcrq1 mega_shift_0_reg_2__15_ ( .D(N870), .SD(mega_shift_0[46]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[47]) );
  sdcrq1 mega_shift_0_reg_1__15_ ( .D(N630), .SD(mega_shift_0[62]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[63]) );
  sdcfq1 mega_shift_1_reg_4__15_ ( .D(sd_wfifo_DQ_in[31]), .SD(
        mega_shift_1_14_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), 
        .Q(test_so2) );
  sdcfq1 mega_shift_1_reg_3__15_ ( .D(N2070), .SD(mega_shift_1_30_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_31_) );
  sdcfq1 mega_shift_1_reg_2__15_ ( .D(N1830), .SD(mega_shift_1_46_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_47_) );
  sdcfq1 mega_shift_1_reg_1__15_ ( .D(N1590), .SD(mega_shift_1_62_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_63_) );
  sdcrq1 mega_shift_0_reg_4__11_ ( .D(sd_wfifo_DQ_in[11]), .SD(
        mega_shift_0[10]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_0[11]) );
  sdcrq1 mega_shift_0_reg_4__5_ ( .D(sd_wfifo_DQ_in[5]), .SD(mega_shift_0[4]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[5])
         );
  sdcrq1 mega_shift_0_reg_4__1_ ( .D(sd_wfifo_DQ_in[1]), .SD(mega_shift_0[0]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[1])
         );
  sdcrq1 mega_shift_0_reg_3__5_ ( .D(N990), .SD(mega_shift_0[20]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[21]) );
  sdcrq1 mega_shift_0_reg_3__1_ ( .D(N990), .SD(mega_shift_0[16]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[17]) );
  sdcrq1 mega_shift_0_reg_3__11_ ( .D(N990), .SD(mega_shift_0[26]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[27]) );
  sdcrq1 mega_shift_0_reg_2__11_ ( .D(N870), .SD(mega_shift_0[42]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[43]) );
  sdcrq1 mega_shift_0_reg_2__5_ ( .D(N870), .SD(mega_shift_0[36]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[37]) );
  sdcrq1 mega_shift_0_reg_2__1_ ( .D(N870), .SD(mega_shift_0[32]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[33]) );
  sdcrq1 mega_shift_0_reg_1__11_ ( .D(N630), .SD(mega_shift_0[58]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[59]) );
  sdcrq1 mega_shift_0_reg_1__5_ ( .D(N630), .SD(mega_shift_0[52]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[53]) );
  sdcrq1 mega_shift_0_reg_1__1_ ( .D(N630), .SD(mega_shift_0[48]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[49]) );
  sdcfq1 mega_shift_1_reg_4__11_ ( .D(sd_wfifo_DQ_in[27]), .SD(
        mega_shift_1_10_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_1_11_) );
  sdcfq1 mega_shift_1_reg_4__5_ ( .D(sd_wfifo_DQ_in[21]), .SD(mega_shift_1_4_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_5_)
         );
  sdcfq1 mega_shift_1_reg_4__1_ ( .D(sd_wfifo_DQ_in[17]), .SD(mega_shift_1_0_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_1_)
         );
  sdcfq1 mega_shift_1_reg_3__11_ ( .D(N2070), .SD(mega_shift_1_26_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_27_) );
  sdcfq1 mega_shift_1_reg_3__5_ ( .D(N2070), .SD(mega_shift_1_20_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_21_) );
  sdcfq1 mega_shift_1_reg_3__1_ ( .D(N2070), .SD(mega_shift_1_16_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_17_) );
  sdcfq1 mega_shift_1_reg_2__11_ ( .D(N1830), .SD(mega_shift_1_42_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_43_) );
  sdcfq1 mega_shift_1_reg_2__5_ ( .D(N1830), .SD(mega_shift_1_36_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_37_) );
  sdcfq1 mega_shift_1_reg_2__1_ ( .D(N1830), .SD(mega_shift_1_32_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_33_) );
  sdcfq1 mega_shift_1_reg_1__11_ ( .D(N1590), .SD(mega_shift_1_58_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_59_) );
  sdcfq1 mega_shift_1_reg_1__5_ ( .D(N1590), .SD(mega_shift_1_52_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_53_) );
  sdcfq1 mega_shift_1_reg_1__1_ ( .D(N1590), .SD(mega_shift_1_48_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_49_) );
  sdcrq1 mega_shift_0_reg_4__8_ ( .D(sd_wfifo_DQ_in[8]), .SD(mega_shift_0[7]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[8])
         );
  sdcrq1 mega_shift_0_reg_4__6_ ( .D(sd_wfifo_DQ_in[6]), .SD(mega_shift_0[5]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[6])
         );
  sdcrq1 mega_shift_0_reg_4__2_ ( .D(sd_wfifo_DQ_in[2]), .SD(mega_shift_0[1]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[2])
         );
  sdcrq1 mega_shift_0_reg_3__8_ ( .D(N990), .SD(mega_shift_0[23]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[24]) );
  sdcrq1 mega_shift_0_reg_3__2_ ( .D(N990), .SD(mega_shift_0[17]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[18]) );
  sdcrq1 mega_shift_0_reg_3__6_ ( .D(N990), .SD(mega_shift_0[21]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[22]) );
  sdcrq1 mega_shift_0_reg_2__2_ ( .D(N870), .SD(mega_shift_0[33]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[34]) );
  sdcrq1 mega_shift_0_reg_2__6_ ( .D(N870), .SD(mega_shift_0[37]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[38]) );
  sdcrq1 mega_shift_0_reg_2__8_ ( .D(N870), .SD(mega_shift_0[39]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[40]) );
  sdcrq1 mega_shift_0_reg_1__2_ ( .D(N630), .SD(mega_shift_0[49]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[50]) );
  sdcrq1 mega_shift_0_reg_1__6_ ( .D(N630), .SD(mega_shift_0[53]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[54]) );
  sdcrq1 mega_shift_0_reg_1__8_ ( .D(N630), .SD(mega_shift_0[55]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[56]) );
  sdcfq1 mega_shift_1_reg_4__8_ ( .D(sd_wfifo_DQ_in[24]), .SD(mega_shift_1_7_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_8_)
         );
  sdcfq1 mega_shift_1_reg_4__6_ ( .D(sd_wfifo_DQ_in[22]), .SD(mega_shift_1_5_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_6_)
         );
  sdcfq1 mega_shift_1_reg_4__2_ ( .D(sd_wfifo_DQ_in[18]), .SD(mega_shift_1_1_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_2_)
         );
  sdcfq1 mega_shift_1_reg_3__2_ ( .D(N2070), .SD(mega_shift_1_17_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_18_) );
  sdcfq1 mega_shift_1_reg_3__6_ ( .D(N2070), .SD(mega_shift_1_21_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_22_) );
  sdcfq1 mega_shift_1_reg_3__8_ ( .D(N2070), .SD(mega_shift_1_23_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_24_) );
  sdcfq1 mega_shift_1_reg_2__2_ ( .D(N1830), .SD(mega_shift_1_33_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_34_) );
  sdcfq1 mega_shift_1_reg_2__6_ ( .D(N1830), .SD(mega_shift_1_37_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_38_) );
  sdcfq1 mega_shift_1_reg_2__8_ ( .D(N1830), .SD(mega_shift_1_39_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_40_) );
  sdcfq1 mega_shift_1_reg_1__2_ ( .D(N1590), .SD(mega_shift_1_49_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_50_) );
  sdcfq1 mega_shift_1_reg_1__6_ ( .D(N1590), .SD(mega_shift_1_53_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_54_) );
  sdcfq1 mega_shift_1_reg_1__8_ ( .D(N1590), .SD(mega_shift_1_55_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_56_) );
  sdcrq1 mega_shift_0_reg_4__9_ ( .D(sd_wfifo_DQ_in[9]), .SD(mega_shift_0[8]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[9])
         );
  sdcrq1 mega_shift_0_reg_4__7_ ( .D(sd_wfifo_DQ_in[7]), .SD(mega_shift_0[6]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[7])
         );
  sdcrq1 mega_shift_0_reg_4__3_ ( .D(sd_wfifo_DQ_in[3]), .SD(mega_shift_0[2]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[3])
         );
  sdcrq1 mega_shift_0_reg_3__7_ ( .D(N990), .SD(mega_shift_0[22]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[23]) );
  sdcrq1 mega_shift_0_reg_3__3_ ( .D(N990), .SD(mega_shift_0[18]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[19]) );
  sdcrq1 mega_shift_0_reg_3__9_ ( .D(N990), .SD(mega_shift_0[24]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[25]) );
  sdcrq1 mega_shift_0_reg_2__9_ ( .D(N870), .SD(mega_shift_0[40]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[41]) );
  sdcrq1 mega_shift_0_reg_2__7_ ( .D(N870), .SD(mega_shift_0[38]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[39]) );
  sdcrq1 mega_shift_0_reg_2__3_ ( .D(N870), .SD(mega_shift_0[34]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[35]) );
  sdcrq1 mega_shift_0_reg_1__9_ ( .D(N630), .SD(mega_shift_0[56]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[57]) );
  sdcrq1 mega_shift_0_reg_1__7_ ( .D(N630), .SD(mega_shift_0[54]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[55]) );
  sdcrq1 mega_shift_0_reg_1__3_ ( .D(N630), .SD(mega_shift_0[50]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[51]) );
  sdcfq1 mega_shift_1_reg_4__9_ ( .D(sd_wfifo_DQ_in[25]), .SD(mega_shift_1_8_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_9_)
         );
  sdcfq1 mega_shift_1_reg_4__7_ ( .D(sd_wfifo_DQ_in[23]), .SD(mega_shift_1_6_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_7_)
         );
  sdcfq1 mega_shift_1_reg_4__3_ ( .D(sd_wfifo_DQ_in[19]), .SD(mega_shift_1_2_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_3_)
         );
  sdcfq1 mega_shift_1_reg_3__9_ ( .D(N2070), .SD(mega_shift_1_24_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_25_) );
  sdcfq1 mega_shift_1_reg_3__7_ ( .D(N2070), .SD(mega_shift_1_22_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_23_) );
  sdcfq1 mega_shift_1_reg_3__3_ ( .D(N2070), .SD(mega_shift_1_18_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_19_) );
  sdcfq1 mega_shift_1_reg_2__9_ ( .D(N1830), .SD(mega_shift_1_40_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_41_) );
  sdcfq1 mega_shift_1_reg_2__7_ ( .D(N1830), .SD(mega_shift_1_38_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_39_) );
  sdcfq1 mega_shift_1_reg_2__3_ ( .D(N1830), .SD(mega_shift_1_34_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_35_) );
  sdcfq1 mega_shift_1_reg_1__9_ ( .D(N1590), .SD(mega_shift_1_56_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_57_) );
  sdcfq1 mega_shift_1_reg_1__7_ ( .D(N1590), .SD(mega_shift_1_54_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_55_) );
  sdcfq1 mega_shift_1_reg_1__3_ ( .D(N1590), .SD(mega_shift_1_50_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_51_) );
  sdcrq1 mega_shift_0_reg_4__14_ ( .D(sd_wfifo_DQ_in[14]), .SD(
        mega_shift_0[13]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_0[14]) );
  sdcrq1 mega_shift_0_reg_4__13_ ( .D(sd_wfifo_DQ_in[13]), .SD(
        mega_shift_0[12]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_0[13]) );
  sdcrq1 mega_shift_0_reg_4__10_ ( .D(sd_wfifo_DQ_in[10]), .SD(mega_shift_0[9]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[10]) );
  sdcrq1 mega_shift_0_reg_4__4_ ( .D(sd_wfifo_DQ_in[4]), .SD(mega_shift_0[3]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[4])
         );
  sdcrq1 mega_shift_0_reg_4__0_ ( .D(sd_wfifo_DQ_in[0]), .SD(mega_shift_0[31]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[0])
         );
  sdcrq1 mega_shift_0_reg_3__13_ ( .D(N990), .SD(mega_shift_0[28]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[29]) );
  sdcrq1 mega_shift_0_reg_3__10_ ( .D(N990), .SD(mega_shift_0[25]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[26]) );
  sdcrq1 mega_shift_0_reg_3__14_ ( .D(N990), .SD(mega_shift_0[29]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[30]) );
  sdcrq1 mega_shift_0_reg_3__0_ ( .D(N990), .SD(mega_shift_0[47]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[16]) );
  sdcrq1 mega_shift_0_reg_3__4_ ( .D(N990), .SD(mega_shift_0[19]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[20]) );
  sdcrq1 mega_shift_0_reg_2__13_ ( .D(N870), .SD(mega_shift_0[44]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[45]) );
  sdcrq1 mega_shift_0_reg_2__0_ ( .D(N870), .SD(mega_shift_0[63]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[32]) );
  sdcrq1 mega_shift_0_reg_2__4_ ( .D(N870), .SD(mega_shift_0[35]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[36]) );
  sdcrq1 mega_shift_0_reg_2__10_ ( .D(N870), .SD(mega_shift_0[41]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[42]) );
  sdcrq1 mega_shift_0_reg_2__14_ ( .D(N870), .SD(mega_shift_0[45]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[46]) );
  sdcrq1 mega_shift_0_reg_1__13_ ( .D(N630), .SD(mega_shift_0[60]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[61]) );
  sdcrq1 mega_shift_0_reg_1__0_ ( .D(N630), .SD(mega_shift_0[79]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[48]) );
  sdcrq1 mega_shift_0_reg_1__4_ ( .D(N630), .SD(mega_shift_0[51]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[52]) );
  sdcrq1 mega_shift_0_reg_1__10_ ( .D(N630), .SD(mega_shift_0[57]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[58]) );
  sdcrq1 mega_shift_0_reg_1__14_ ( .D(N630), .SD(mega_shift_0[61]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[62]) );
  sdcfq1 mega_shift_1_reg_4__14_ ( .D(sd_wfifo_DQ_in[30]), .SD(
        mega_shift_1_13_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_1_14_) );
  sdcfq1 mega_shift_1_reg_4__13_ ( .D(sd_wfifo_DQ_in[29]), .SD(
        mega_shift_1_12_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_1_13_) );
  sdcfq1 mega_shift_1_reg_4__10_ ( .D(sd_wfifo_DQ_in[26]), .SD(mega_shift_1_9_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_10_) );
  sdcfq1 mega_shift_1_reg_4__4_ ( .D(sd_wfifo_DQ_in[20]), .SD(mega_shift_1_3_), 
        .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_4_)
         );
  sdcfq1 mega_shift_1_reg_4__0_ ( .D(sd_wfifo_DQ_in[16]), .SD(mega_shift_1_31_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_0_) );
  sdcfq1 mega_shift_1_reg_3__13_ ( .D(N2070), .SD(mega_shift_1_28_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_29_) );
  sdcfq1 mega_shift_1_reg_3__0_ ( .D(N2070), .SD(mega_shift_1_47_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_16_) );
  sdcfq1 mega_shift_1_reg_3__4_ ( .D(N2070), .SD(mega_shift_1_19_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_20_) );
  sdcfq1 mega_shift_1_reg_3__10_ ( .D(N2070), .SD(mega_shift_1_25_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_26_) );
  sdcfq1 mega_shift_1_reg_3__14_ ( .D(N2070), .SD(mega_shift_1_29_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_30_) );
  sdcfq1 mega_shift_1_reg_2__13_ ( .D(N1830), .SD(mega_shift_1_44_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_45_) );
  sdcfq1 mega_shift_1_reg_2__0_ ( .D(N1830), .SD(mega_shift_1_63_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_32_) );
  sdcfq1 mega_shift_1_reg_2__4_ ( .D(N1830), .SD(mega_shift_1_35_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_36_) );
  sdcfq1 mega_shift_1_reg_2__10_ ( .D(N1830), .SD(mega_shift_1_41_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_42_) );
  sdcfq1 mega_shift_1_reg_2__14_ ( .D(N1830), .SD(mega_shift_1_45_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_46_) );
  sdcfq1 mega_shift_1_reg_1__13_ ( .D(N1590), .SD(mega_shift_1_60_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_61_) );
  sdcfq1 mega_shift_1_reg_1__0_ ( .D(N1590), .SD(mega_shift_1_79_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_48_) );
  sdcfq1 mega_shift_1_reg_1__4_ ( .D(N1590), .SD(mega_shift_1_51_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_52_) );
  sdcfq1 mega_shift_1_reg_1__10_ ( .D(N1590), .SD(mega_shift_1_57_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_58_) );
  sdcfq1 mega_shift_1_reg_1__14_ ( .D(N1590), .SD(mega_shift_1_61_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_62_) );
  sdcrq1 mega_shift_0_reg_4__12_ ( .D(sd_wfifo_DQ_in[12]), .SD(
        mega_shift_0[11]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_0[12]) );
  sdcrq1 mega_shift_0_reg_3__12_ ( .D(N990), .SD(mega_shift_0[27]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[28]) );
  sdcrq1 mega_shift_0_reg_2__12_ ( .D(N870), .SD(mega_shift_0[43]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[44]) );
  sdcrq1 mega_shift_0_reg_1__12_ ( .D(N630), .SD(mega_shift_0[59]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[60]) );
  sdcfq1 mega_shift_1_reg_4__12_ ( .D(sd_wfifo_DQ_in[28]), .SD(
        mega_shift_1_11_), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), 
        .Q(mega_shift_1_12_) );
  sdcfq1 mega_shift_1_reg_3__12_ ( .D(N2070), .SD(mega_shift_1_27_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_28_) );
  sdcfq1 mega_shift_1_reg_2__12_ ( .D(N1830), .SD(mega_shift_1_43_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_44_) );
  sdcfq1 mega_shift_1_reg_1__12_ ( .D(N1590), .SD(mega_shift_1_59_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_60_) );
  sdnrq1 control_bus_reg_14_ ( .D(test_so1), .SD(n321), .SC(test_se), .CP(
        sdram_clk), .Q(control_bus[14]) );
  sdnrq1 control_bus_reg_7_ ( .D(sync_control_bus_7_), .SD(n473), .SC(test_se), 
        .CP(sdram_clk), .Q(control_bus[7]) );
  sdcrq1 out_control_reg_14_ ( .D(c_out_control[14]), .SD(sd_BWS[0]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_wfifo_pop) );
  sdnrq1 control_bus_reg_10_ ( .D(sync_control_bus_10_), .SD(control_bus[9]), 
        .SC(test_se), .CP(sdram_clk), .Q(control_bus[10]) );
  sdnrq1 control_bus_reg_6_ ( .D(sync_control_bus_6_), .SD(control_bus[5]), 
        .SC(test_se), .CP(sdram_clk), .Q(control_bus[6]) );
  sdnrq1 control_bus_reg_2_ ( .D(sync_control_bus_2_), .SD(n371), .SC(test_se), 
        .CP(sdram_clk), .Q(add_155_carry_6_) );
  sdcrq1 out_control_reg_15_ ( .D(c_out_control[15]), .SD(sd_wfifo_pop), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_rfifo_push) );
  sdnrq1 control_bus_reg_9_ ( .D(sync_control_bus_9_), .SD(control_bus[8]), 
        .SC(test_se), .CP(sdram_clk), .Q(control_bus[9]) );
  sdnrq1 control_bus_reg_4_ ( .D(sync_control_bus_4_), .SD(control_bus[3]), 
        .SC(test_se), .CP(sdram_clk), .Q(control_bus[4]) );
  sdnrq1 control_bus_reg_5_ ( .D(sync_control_bus_5_), .SD(control_bus[4]), 
        .SC(test_se), .CP(sdram_clk), .Q(control_bus[5]) );
  sdnrq1 control_bus_reg_0_ ( .D(sync_control_bus_0_), .SD(DQ_out_0[15]), .SC(
        test_se), .CP(sdram_clk), .Q(N41) );
  sdnrq1 control_bus_reg_1_ ( .D(sync_control_bus_1_), .SD(n363), .SC(test_se), 
        .CP(sdram_clk), .Q(N42) );
  sdnrq1 sync_control_bus_reg_6_ ( .D(risc_PSW[2]), .SD(sync_control_bus_5_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_6_) );
  sdnrq1 sync_control_bus_reg_5_ ( .D(risc_PSW[1]), .SD(sync_control_bus_4_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_5_) );
  sdnrq1 sync_control_bus_reg_4_ ( .D(risc_PSW[0]), .SD(sync_control_bus_3_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_4_) );
  sdcrq1 mega_shift_0_reg_0__15_ ( .D(N390), .SD(mega_shift_0[78]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[79]) );
  sdcrq1 mega_shift_0_reg_0__13_ ( .D(N390), .SD(mega_shift_0[76]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[77]) );
  sdcrq1 mega_shift_0_reg_0__11_ ( .D(N390), .SD(mega_shift_0[74]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[75]) );
  sdcrq1 mega_shift_0_reg_0__9_ ( .D(N390), .SD(mega_shift_0[72]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[73]) );
  sdcrq1 mega_shift_0_reg_0__7_ ( .D(N390), .SD(mega_shift_0[70]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[71]) );
  sdcrq1 mega_shift_0_reg_0__5_ ( .D(N390), .SD(mega_shift_0[68]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[69]) );
  sdcrq1 mega_shift_0_reg_0__3_ ( .D(N390), .SD(mega_shift_0[66]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[67]) );
  sdcrq1 mega_shift_0_reg_0__1_ ( .D(N390), .SD(mega_shift_0[64]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[65]) );
  sdcrq1 mega_shift_0_reg_0__0_ ( .D(N390), .SD(control_bus[14]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[64]) );
  sdcrq1 mega_shift_0_reg_0__2_ ( .D(N390), .SD(mega_shift_0[65]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[66]) );
  sdcrq1 mega_shift_0_reg_0__4_ ( .D(N390), .SD(mega_shift_0[67]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[68]) );
  sdcrq1 mega_shift_0_reg_0__6_ ( .D(N390), .SD(mega_shift_0[69]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[70]) );
  sdcrq1 mega_shift_0_reg_0__8_ ( .D(N390), .SD(mega_shift_0[71]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[72]) );
  sdcrq1 mega_shift_0_reg_0__10_ ( .D(N390), .SD(mega_shift_0[73]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[74]) );
  sdcrq1 mega_shift_0_reg_0__12_ ( .D(N390), .SD(mega_shift_0[75]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[76]) );
  sdcrq1 mega_shift_0_reg_0__14_ ( .D(N390), .SD(mega_shift_0[77]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_0[78]) );
  sdcfq1 mega_shift_1_reg_0__15_ ( .D(N1350), .SD(mega_shift_1_78_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_79_) );
  sdcfq1 mega_shift_1_reg_0__13_ ( .D(N1350), .SD(mega_shift_1_76_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_77_) );
  sdcfq1 mega_shift_1_reg_0__11_ ( .D(N1350), .SD(mega_shift_1_74_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_75_) );
  sdcfq1 mega_shift_1_reg_0__9_ ( .D(N1350), .SD(mega_shift_1_72_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_73_) );
  sdcfq1 mega_shift_1_reg_0__7_ ( .D(N1350), .SD(mega_shift_1_70_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_71_) );
  sdcfq1 mega_shift_1_reg_0__5_ ( .D(N1350), .SD(mega_shift_1_68_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_69_) );
  sdcfq1 mega_shift_1_reg_0__3_ ( .D(N1350), .SD(mega_shift_1_66_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_67_) );
  sdcfq1 mega_shift_1_reg_0__1_ ( .D(N1350), .SD(mega_shift_1_64_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_65_) );
  sdcfq1 mega_shift_1_reg_0__0_ ( .D(N1350), .SD(DQ_out_1[15]), .SC(test_se), 
        .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_64_) );
  sdcfq1 mega_shift_1_reg_0__2_ ( .D(N1350), .SD(mega_shift_1_65_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_66_) );
  sdcfq1 mega_shift_1_reg_0__4_ ( .D(N1350), .SD(mega_shift_1_67_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_68_) );
  sdcfq1 mega_shift_1_reg_0__6_ ( .D(N1350), .SD(mega_shift_1_69_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_70_) );
  sdcfq1 mega_shift_1_reg_0__8_ ( .D(N1350), .SD(mega_shift_1_71_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_72_) );
  sdcfq1 mega_shift_1_reg_0__10_ ( .D(N1350), .SD(mega_shift_1_73_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_74_) );
  sdcfq1 mega_shift_1_reg_0__12_ ( .D(N1350), .SD(mega_shift_1_75_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_76_) );
  sdcfq1 mega_shift_1_reg_0__14_ ( .D(N1350), .SD(mega_shift_1_77_), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(mega_shift_1_78_) );
  sdcrq1 out_control_reg_12_ ( .D(c_out_control[12]), .SD(sd_RW), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_BWS[0]) );
  sdcrq1 out_control_reg_8_ ( .D(c_out_control[8]), .SD(sd_A[7]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[8]) );
  sdcrq1 out_control_reg_7_ ( .D(c_out_control[7]), .SD(sd_A[6]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[7]) );
  sdcrq1 out_control_reg_4_ ( .D(c_out_control[4]), .SD(sd_A[3]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[4]) );
  sdnrq1 sync_control_bus_reg_3_ ( .D(risc_OUT_VALID), .SD(sync_control_bus_2_), .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_3_) );
  sdnrq1 sync_control_bus_reg_0_ ( .D(risc_Rd_Instr), .SD(sd_DQ_en[15]), .SC(
        test_se), .CP(sdram_clk), .Q(sync_control_bus_0_) );
  sdcrq1 out_control_reg_13_ ( .D(c_out_control[13]), .SD(test_si3), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_BWS[1]) );
  sdcrq1 out_control_reg_11_ ( .D(c_out_control[11]), .SD(sd_LD), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_RW) );
  sdcrq1 out_control_reg_9_ ( .D(c_out_control[9]), .SD(sd_A[8]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[9]) );
  sdcrq1 out_control_reg_6_ ( .D(c_out_control[6]), .SD(sd_A[5]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[6]) );
  sdcrq1 out_control_reg_3_ ( .D(c_out_control[3]), .SD(sd_A[2]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[3]) );
  sdcrq1 out_control_reg_2_ ( .D(c_out_control[2]), .SD(sd_A[1]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[2]) );
  sdcrq1 out_control_reg_10_ ( .D(c_out_control[10]), .SD(sd_A[9]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_LD) );
  sdcrq1 out_control_reg_5_ ( .D(c_out_control[5]), .SD(sd_A[4]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[5]) );
  sdcrq1 out_control_reg_1_ ( .D(c_out_control[1]), .SD(sd_A[0]), .SC(test_se), 
        .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[1]) );
  sdcrq1 out_control_reg_0_ ( .D(c_out_control[0]), .SD(mega_shift_0[15]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(sd_A[0]) );
  sdnrq1 sync_control_bus_reg_14_ ( .D(risc_PSW[10]), .SD(sync_control_bus_13_), .SC(test_se), .CP(sdram_clk), .Q(test_so1) );
  sdnrq1 sync_control_bus_reg_13_ ( .D(risc_PSW[9]), .SD(sync_control_bus_12_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_13_) );
  sdnrq1 sync_control_bus_reg_12_ ( .D(risc_PSW[8]), .SD(sync_control_bus_11_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_12_) );
  sdnrq1 sync_control_bus_reg_11_ ( .D(risc_PSW[7]), .SD(sync_control_bus_10_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_11_) );
  sdnrq1 sync_control_bus_reg_10_ ( .D(risc_PSW[6]), .SD(sync_control_bus_9_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_10_) );
  sdnrq1 sync_control_bus_reg_9_ ( .D(risc_PSW[5]), .SD(sync_control_bus_8_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_9_) );
  sdnrq1 sync_control_bus_reg_8_ ( .D(risc_PSW[4]), .SD(sync_control_bus_7_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_8_) );
  sdnrq1 sync_control_bus_reg_7_ ( .D(risc_PSW[3]), .SD(sync_control_bus_6_), 
        .SC(test_se), .CP(sdram_clk), .Q(sync_control_bus_7_) );
  sdnrq1 sync_control_bus_reg_2_ ( .D(risc_STACK_FULL), .SD(
        sync_control_bus_1_), .SC(test_se), .CP(sdram_clk), .Q(
        sync_control_bus_2_) );
  sdnrq1 sync_control_bus_reg_1_ ( .D(risc_EndOfInstrn), .SD(
        sync_control_bus_0_), .SC(test_se), .CP(sdram_clk), .Q(
        sync_control_bus_1_) );
  sdcrq1 DQ_out_0_reg_15_ ( .D(mega_shift_0[79]), .SD(DQ_out_0[14]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[15]) );
  sdcrq1 DQ_out_0_reg_13_ ( .D(mega_shift_0[77]), .SD(DQ_out_0[12]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[13]) );
  sdcrq1 DQ_out_0_reg_11_ ( .D(mega_shift_0[75]), .SD(DQ_out_0[10]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[11]) );
  sdcrq1 DQ_out_0_reg_9_ ( .D(mega_shift_0[73]), .SD(DQ_out_0[8]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[9]) );
  sdcrq1 DQ_out_0_reg_7_ ( .D(mega_shift_0[71]), .SD(DQ_out_0[6]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[7]) );
  sdcrq1 DQ_out_0_reg_5_ ( .D(mega_shift_0[69]), .SD(DQ_out_0[4]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[5]) );
  sdcrq1 DQ_out_0_reg_3_ ( .D(mega_shift_0[67]), .SD(DQ_out_0[2]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[3]) );
  sdcrq1 DQ_out_0_reg_1_ ( .D(mega_shift_0[65]), .SD(DQ_out_0[0]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[1]) );
  sdcrq1 DQ_out_0_reg_0_ ( .D(mega_shift_0[64]), .SD(sd_rfifo_DQ_out[15]), 
        .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[0]) );
  sdcrq1 DQ_out_0_reg_2_ ( .D(mega_shift_0[66]), .SD(DQ_out_0[1]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[2]) );
  sdcrq1 DQ_out_0_reg_4_ ( .D(mega_shift_0[68]), .SD(DQ_out_0[3]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[4]) );
  sdcrq1 DQ_out_0_reg_6_ ( .D(mega_shift_0[70]), .SD(DQ_out_0[5]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[6]) );
  sdcrq1 DQ_out_0_reg_8_ ( .D(mega_shift_0[72]), .SD(DQ_out_0[7]), .SC(test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[8]) );
  sdcrq1 DQ_out_0_reg_10_ ( .D(mega_shift_0[74]), .SD(DQ_out_0[9]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[10]) );
  sdcrq1 DQ_out_0_reg_12_ ( .D(mega_shift_0[76]), .SD(DQ_out_0[11]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[12]) );
  sdcrq1 DQ_out_0_reg_14_ ( .D(mega_shift_0[78]), .SD(DQ_out_0[13]), .SC(
        test_se), .CP(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_0[14]) );
  sdcfq1 DQ_out_1_reg_15_ ( .D(mega_shift_1_79_), .SD(DQ_out_1[14]), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[15]) );
  sdcfq1 DQ_out_1_reg_13_ ( .D(mega_shift_1_77_), .SD(DQ_out_1[12]), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[13]) );
  sdcfq1 DQ_out_1_reg_11_ ( .D(mega_shift_1_75_), .SD(DQ_out_1[10]), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[11]) );
  sdcfq1 DQ_out_1_reg_9_ ( .D(mega_shift_1_73_), .SD(DQ_out_1[8]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[9]) );
  sdcfq1 DQ_out_1_reg_7_ ( .D(mega_shift_1_71_), .SD(DQ_out_1[6]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[7]) );
  sdcfq1 DQ_out_1_reg_5_ ( .D(mega_shift_1_69_), .SD(DQ_out_1[4]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[5]) );
  sdcfq1 DQ_out_1_reg_3_ ( .D(mega_shift_1_67_), .SD(DQ_out_1[2]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[3]) );
  sdcfq1 DQ_out_1_reg_1_ ( .D(mega_shift_1_65_), .SD(DQ_out_1[0]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[1]) );
  sdcfq1 DQ_out_1_reg_0_ ( .D(mega_shift_1_64_), .SD(n503), .SC(test_se), 
        .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[0]) );
  sdcfq1 DQ_out_1_reg_2_ ( .D(mega_shift_1_66_), .SD(DQ_out_1[1]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[2]) );
  sdcfq1 DQ_out_1_reg_4_ ( .D(mega_shift_1_68_), .SD(DQ_out_1[3]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[4]) );
  sdcfq1 DQ_out_1_reg_6_ ( .D(mega_shift_1_70_), .SD(DQ_out_1[5]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[6]) );
  sdcfq1 DQ_out_1_reg_8_ ( .D(mega_shift_1_72_), .SD(DQ_out_1[7]), .SC(test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[8]) );
  sdcfq1 DQ_out_1_reg_10_ ( .D(mega_shift_1_74_), .SD(DQ_out_1[9]), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[10]) );
  sdcfq1 DQ_out_1_reg_12_ ( .D(mega_shift_1_76_), .SD(DQ_out_1[11]), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[12]) );
  sdcfq1 DQ_out_1_reg_14_ ( .D(mega_shift_1_78_), .SD(DQ_out_1[13]), .SC(
        test_se), .CPN(sdram_clk), .CDN(sdram_rst_n), .Q(DQ_out_1[14]) );
  sdcrq1 sd_DQ_en_reg_0_ ( .D(N7), .SD(sd_rfifo_push), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n499) );
  sdcrq1 sd_DQ_en_reg_1_ ( .D(N7), .SD(sd_DQ_en[0]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n498) );
  sdcrq1 sd_DQ_en_reg_2_ ( .D(N7), .SD(sd_DQ_en[1]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n497) );
  sdcrq1 sd_DQ_en_reg_3_ ( .D(N7), .SD(sd_DQ_en[2]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n496) );
  sdcrq1 sd_DQ_en_reg_4_ ( .D(N7), .SD(sd_DQ_en[3]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n495) );
  sdcrq1 sd_DQ_en_reg_5_ ( .D(N7), .SD(sd_DQ_en[4]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n494) );
  sdcrq1 sd_DQ_en_reg_6_ ( .D(N7), .SD(sd_DQ_en[5]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n493) );
  sdcrq1 sd_DQ_en_reg_7_ ( .D(N7), .SD(sd_DQ_en[6]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n492) );
  sdcrq1 sd_DQ_en_reg_8_ ( .D(N7), .SD(sd_DQ_en[7]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n491) );
  sdcrq1 sd_DQ_en_reg_9_ ( .D(N7), .SD(sd_DQ_en[8]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n490) );
  sdcrq1 sd_DQ_en_reg_15_ ( .D(N7), .SD(sd_DQ_en[14]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n484) );
  sdcrq1 sd_DQ_en_reg_10_ ( .D(N7), .SD(sd_DQ_en[9]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n489) );
  sdcrq1 sd_DQ_en_reg_14_ ( .D(N7), .SD(sd_DQ_en[13]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n485) );
  sdcrq1 sd_DQ_en_reg_11_ ( .D(N7), .SD(sd_DQ_en[10]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n488) );
  sdcrq1 sd_DQ_en_reg_13_ ( .D(N7), .SD(sd_DQ_en[12]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n486) );
  sdcrq1 sd_DQ_en_reg_12_ ( .D(N7), .SD(sd_DQ_en[11]), .SC(test_se), .CP(
        sdram_clk), .CDN(sdram_rst_n), .Q(n487) );
  bufbd7 U5 ( .I(n487), .Z(sd_DQ_en[12]) );
  bufbd7 U6 ( .I(n486), .Z(sd_DQ_en[13]) );
  bufbd7 U7 ( .I(n488), .Z(sd_DQ_en[11]) );
  bufbd7 U8 ( .I(n485), .Z(sd_DQ_en[14]) );
  bufbd7 U9 ( .I(n489), .Z(sd_DQ_en[10]) );
  bufbd7 U10 ( .I(n484), .Z(sd_DQ_en[15]) );
  bufbd7 U11 ( .I(n490), .Z(sd_DQ_en[9]) );
  bufbd7 U12 ( .I(n491), .Z(sd_DQ_en[8]) );
  bufbd7 U274 ( .I(n492), .Z(sd_DQ_en[7]) );
  bufbd7 U285 ( .I(n493), .Z(sd_DQ_en[6]) );
  bufbd7 U292 ( .I(n494), .Z(sd_DQ_en[5]) );
  bufbd7 U295 ( .I(n495), .Z(sd_DQ_en[4]) );
  bufbd7 U298 ( .I(n496), .Z(sd_DQ_en[3]) );
  bufbd7 U302 ( .I(n497), .Z(sd_DQ_en[2]) );
  bufbd7 U303 ( .I(n498), .Z(sd_DQ_en[1]) );
  bufbd7 U304 ( .I(n499), .Z(sd_DQ_en[0]) );
  inv0d1 U305 ( .I(c_out_control[0]), .ZN(N7) );
  bufbd1 U306 ( .I(sd_wfifo_empty), .Z(n483) );
  inv0d1 U307 ( .I(n367), .ZN(n328) );
  nd12d0 U308 ( .A1(n333), .A2(n364), .ZN(c_out_control[0]) );
  nd02d1 U309 ( .A1(n349), .A2(n350), .ZN(c_out_control[1]) );
  nd02d1 U310 ( .A1(n341), .A2(n342), .ZN(c_out_control[5]) );
  nd02d1 U311 ( .A1(n361), .A2(n362), .ZN(c_out_control[10]) );
  inv0d1 U312 ( .I(n365), .ZN(n330) );
  nd02d1 U313 ( .A1(n359), .A2(n360), .ZN(c_out_control[11]) );
  nd02d1 U314 ( .A1(n355), .A2(n356), .ZN(c_out_control[13]) );
  nd02d1 U315 ( .A1(n353), .A2(n354), .ZN(c_out_control[14]) );
  nd02d1 U316 ( .A1(n351), .A2(n352), .ZN(c_out_control[15]) );
  inv0d1 U317 ( .I(n17), .ZN(n372) );
  inv0d1 U318 ( .I(n17), .ZN(n383) );
  inv0d1 U319 ( .I(n17), .ZN(n363) );
  an03d1 U320 ( .A1(n388), .A2(n389), .A3(n375), .Z(n333) );
  an04d1 U321 ( .A1(n375), .A2(n388), .A3(n374), .A4(n387), .Z(n331) );
  an04d1 U322 ( .A1(n374), .A2(n373), .A3(n386), .A4(n387), .Z(n334) );
  an04d1 U324 ( .A1(n366), .A2(n365), .A3(n367), .A4(n368), .Z(n327) );
  an03d1 U325 ( .A1(n373), .A2(n386), .A3(n389), .Z(n332) );
  inv0d1 U326 ( .I(control_bus[8]), .ZN(n391) );
  nd02d1 U327 ( .A1(n347), .A2(n348), .ZN(c_out_control[2]) );
  nd02d1 U328 ( .A1(n345), .A2(n346), .ZN(c_out_control[3]) );
  nd02d1 U329 ( .A1(n339), .A2(n340), .ZN(c_out_control[6]) );
  nd02d1 U335 ( .A1(n325), .A2(n326), .ZN(c_out_control[9]) );
  inv0d1 U336 ( .I(n466), .ZN(n468) );
  inv0d1 U337 ( .I(n470), .ZN(n472) );
  inv0d1 U338 ( .I(n466), .ZN(n469) );
  inv0d1 U340 ( .I(n470), .ZN(n473) );
  inv0d1 U341 ( .I(n478), .ZN(n481) );
  inv0d1 U342 ( .I(n470), .ZN(n471) );
  inv0d1 U343 ( .I(n466), .ZN(n467) );
  inv0d1 U344 ( .I(n476), .ZN(n380) );
  inv0d1 U345 ( .I(n366), .ZN(n329) );
  inv0d1 U346 ( .I(n474), .ZN(n476) );
  inv0d1 U347 ( .I(n474), .ZN(n477) );
  inv0d1 U348 ( .I(n478), .ZN(n480) );
  inv0d1 U349 ( .I(control_bus[13]), .ZN(n385) );
  inv0d1 U350 ( .I(n474), .ZN(n475) );
  inv0d1 U351 ( .I(n478), .ZN(n479) );
  bufbd1 U352 ( .I(sd_rfifo_full), .Z(n482) );
  inv0d1 U353 ( .I(N41), .ZN(n17) );
  nd02d1 U354 ( .A1(n357), .A2(n358), .ZN(c_out_control[12]) );
  inv0d1 U355 ( .I(n308), .ZN(control_bus[8]) );
  inv0d1 U356 ( .I(n369), .ZN(n384) );
  inv0d1 U357 ( .I(control_bus[12]), .ZN(n393) );
  inv0d1 U358 ( .I(n318), .ZN(control_bus[12]) );
  inv0d1 U359 ( .I(n297), .ZN(control_bus[3]) );
  inv0d1 U360 ( .I(n315), .ZN(control_bus[11]) );
  inv0d1 U361 ( .I(control_bus[6]), .ZN(n470) );
  inv0d1 U362 ( .I(control_bus[10]), .ZN(n478) );
  inv0d1 U363 ( .I(add_155_carry_6_), .ZN(n466) );
  nd02d1 U364 ( .A1(n343), .A2(n344), .ZN(c_out_control[4]) );
  nd02d1 U365 ( .A1(n337), .A2(n338), .ZN(c_out_control[7]) );
  nd02d1 U366 ( .A1(n335), .A2(n336), .ZN(c_out_control[8]) );
  xr03d1 U367 ( .A1(n448), .A2(n449), .A3(n450), .Z(N1350) );
  xr03d1 U368 ( .A1(mega_shift_1_63_), .A2(mega_shift_1_62_), .A3(n452), .Z(
        n449) );
  xr03d1 U369 ( .A1(mega_shift_1_59_), .A2(mega_shift_1_58_), .A3(n451), .Z(
        n450) );
  xr03d1 U370 ( .A1(n439), .A2(n440), .A3(n441), .Z(N1590) );
  xr03d1 U371 ( .A1(mega_shift_1_47_), .A2(mega_shift_1_46_), .A3(n443), .Z(
        n440) );
  xr03d1 U372 ( .A1(mega_shift_1_43_), .A2(mega_shift_1_42_), .A3(n442), .Z(
        n441) );
  xr03d1 U373 ( .A1(n430), .A2(n431), .A3(n432), .Z(N1830) );
  xr03d1 U374 ( .A1(mega_shift_1_31_), .A2(mega_shift_1_30_), .A3(n434), .Z(
        n431) );
  xr03d1 U375 ( .A1(mega_shift_1_27_), .A2(mega_shift_1_26_), .A3(n433), .Z(
        n432) );
  xr03d1 U376 ( .A1(n412), .A2(n413), .A3(n414), .Z(N2070) );
  xr03d1 U377 ( .A1(test_so2), .A2(mega_shift_1_14_), .A3(n416), .Z(n413) );
  xr03d1 U378 ( .A1(mega_shift_1_11_), .A2(mega_shift_1_10_), .A3(n415), .Z(
        n414) );
  xr03d1 U379 ( .A1(n421), .A2(n422), .A3(n423), .Z(N390) );
  xr03d1 U380 ( .A1(mega_shift_0[63]), .A2(mega_shift_0[62]), .A3(n425), .Z(
        n422) );
  xr03d1 U381 ( .A1(mega_shift_0[59]), .A2(mega_shift_0[58]), .A3(n424), .Z(
        n423) );
  xr03d1 U412 ( .A1(n403), .A2(n404), .A3(n405), .Z(N630) );
  xr03d1 U420 ( .A1(mega_shift_0[47]), .A2(mega_shift_0[46]), .A3(n407), .Z(
        n404) );
  xr03d1 U468 ( .A1(mega_shift_0[43]), .A2(mega_shift_0[42]), .A3(n406), .Z(
        n405) );
  xr03d1 U469 ( .A1(n394), .A2(n395), .A3(n396), .Z(N870) );
  xr03d1 U470 ( .A1(mega_shift_0[31]), .A2(mega_shift_0[30]), .A3(n398), .Z(
        n395) );
  xr03d1 U471 ( .A1(mega_shift_0[27]), .A2(mega_shift_0[26]), .A3(n397), .Z(
        n396) );
  xr03d1 U472 ( .A1(n457), .A2(n458), .A3(n459), .Z(N990) );
  xr03d1 U473 ( .A1(mega_shift_0[15]), .A2(mega_shift_0[14]), .A3(n461), .Z(
        n458) );
  xr03d1 U474 ( .A1(mega_shift_0[11]), .A2(mega_shift_0[10]), .A3(n460), .Z(
        n459) );
  inv0d1 U475 ( .I(control_bus[7]), .ZN(n474) );
  inv0d1 U476 ( .I(N42), .ZN(n371) );
  xr03d1 U477 ( .A1(mega_shift_1_49_), .A2(mega_shift_1_48_), .A3(n455), .Z(
        n454) );
  xr03d1 U478 ( .A1(mega_shift_1_33_), .A2(mega_shift_1_32_), .A3(n446), .Z(
        n445) );
  xr03d1 U479 ( .A1(mega_shift_1_17_), .A2(mega_shift_1_16_), .A3(n437), .Z(
        n436) );
  xr03d1 U480 ( .A1(mega_shift_1_1_), .A2(mega_shift_1_0_), .A3(n419), .Z(n418) );
  xr03d1 U481 ( .A1(mega_shift_0[49]), .A2(mega_shift_0[48]), .A3(n428), .Z(
        n427) );
  xr03d1 U482 ( .A1(mega_shift_0[33]), .A2(mega_shift_0[32]), .A3(n410), .Z(
        n409) );
  xr03d1 U483 ( .A1(mega_shift_0[17]), .A2(mega_shift_0[16]), .A3(n401), .Z(
        n400) );
  xr03d1 U484 ( .A1(mega_shift_0[1]), .A2(mega_shift_0[0]), .A3(n464), .Z(n463) );
  inv0d1 U485 ( .I(n321), .ZN(control_bus[13]) );
  xr03d1 U486 ( .A1(mega_shift_1_53_), .A2(mega_shift_1_52_), .A3(n456), .Z(
        n453) );
  xr03d1 U487 ( .A1(mega_shift_1_37_), .A2(mega_shift_1_36_), .A3(n447), .Z(
        n444) );
  xr03d1 U488 ( .A1(mega_shift_1_21_), .A2(mega_shift_1_20_), .A3(n438), .Z(
        n435) );
  xr03d1 U489 ( .A1(mega_shift_1_5_), .A2(mega_shift_1_4_), .A3(n420), .Z(n417) );
  xr03d1 U490 ( .A1(mega_shift_0[53]), .A2(mega_shift_0[52]), .A3(n429), .Z(
        n426) );
  xr03d1 U491 ( .A1(mega_shift_0[37]), .A2(mega_shift_0[36]), .A3(n411), .Z(
        n408) );
  xr03d1 U492 ( .A1(mega_shift_0[21]), .A2(mega_shift_0[20]), .A3(n402), .Z(
        n399) );
  xr03d1 U493 ( .A1(mega_shift_0[5]), .A2(mega_shift_0[4]), .A3(n465), .Z(n462) );
  xr02d1 U494 ( .A1(add_161_carry_15_), .A2(control_bus[12]), .Z(N101) );
  or02d0 U495 ( .A1(add_161_carry_14_), .A2(control_bus[11]), .Z(
        add_161_carry_15_) );
  xn02d1 U496 ( .A1(control_bus[11]), .A2(add_161_carry_14_), .ZN(N100) );
  or02d0 U497 ( .A1(add_161_carry_13_), .A2(n480), .Z(add_161_carry_14_) );
  xn02d1 U498 ( .A1(n480), .A2(add_161_carry_13_), .ZN(N99) );
  an02d0 U499 ( .A1(control_bus[9]), .A2(add_161_carry_12_), .Z(
        add_161_carry_13_) );
  xr02d1 U500 ( .A1(add_161_carry_12_), .A2(control_bus[9]), .Z(N98) );
  or02d0 U501 ( .A1(add_161_carry_11_), .A2(control_bus[8]), .Z(
        add_161_carry_12_) );
  xn02d1 U502 ( .A1(control_bus[8]), .A2(add_161_carry_11_), .ZN(N97) );
  an02d0 U503 ( .A1(n476), .A2(add_161_carry_10_), .Z(add_161_carry_11_) );
  xr02d1 U504 ( .A1(add_161_carry_10_), .A2(n475), .Z(N96) );
  or02d0 U505 ( .A1(add_161_carry_9_), .A2(n471), .Z(add_161_carry_10_) );
  xn02d1 U506 ( .A1(n471), .A2(add_161_carry_9_), .ZN(N95) );
  an02d0 U507 ( .A1(control_bus[5]), .A2(add_161_carry_8_), .Z(
        add_161_carry_9_) );
  xr02d1 U508 ( .A1(add_161_carry_8_), .A2(control_bus[5]), .Z(N94) );
  an02d0 U509 ( .A1(control_bus[4]), .A2(add_161_carry_7_), .Z(
        add_161_carry_8_) );
  xr02d1 U510 ( .A1(add_161_carry_7_), .A2(control_bus[4]), .Z(N93) );
  an02d0 U511 ( .A1(control_bus[3]), .A2(add_161_carry_6_), .Z(
        add_161_carry_7_) );
  xr02d1 U512 ( .A1(add_161_carry_6_), .A2(control_bus[3]), .Z(N92) );
  or02d0 U513 ( .A1(add_161_carry_5_), .A2(n468), .Z(add_161_carry_6_) );
  xn02d1 U514 ( .A1(n468), .A2(add_161_carry_5_), .ZN(N91) );
  or02d0 U515 ( .A1(add_161_carry_4_), .A2(N42), .Z(add_161_carry_5_) );
  xn02d1 U516 ( .A1(N42), .A2(add_161_carry_4_), .ZN(N90) );
  or02d0 U517 ( .A1(add_161_carry_3_), .A2(n372), .Z(add_161_carry_4_) );
  xn02d1 U518 ( .A1(n372), .A2(add_161_carry_3_), .ZN(N89) );
  or02d0 U519 ( .A1(n483), .A2(n482), .Z(add_161_carry_3_) );
  xn02d1 U520 ( .A1(n482), .A2(n483), .ZN(N88) );
  xr02d1 U521 ( .A1(add_163_carry_15_), .A2(control_bus[12]), .Z(N117) );
  or02d0 U522 ( .A1(add_163_carry_14_), .A2(control_bus[11]), .Z(
        add_163_carry_15_) );
  xn02d1 U523 ( .A1(control_bus[11]), .A2(add_163_carry_14_), .ZN(N116) );
  an02d0 U524 ( .A1(n480), .A2(add_163_carry_13_), .Z(add_163_carry_14_) );
  xr02d1 U525 ( .A1(add_163_carry_13_), .A2(n480), .Z(N115) );
  an02d0 U526 ( .A1(control_bus[9]), .A2(add_163_carry_12_), .Z(
        add_163_carry_13_) );
  xr02d1 U527 ( .A1(add_163_carry_12_), .A2(control_bus[9]), .Z(N114) );
  an02d0 U528 ( .A1(control_bus[8]), .A2(add_163_carry_11_), .Z(
        add_163_carry_12_) );
  xr02d1 U529 ( .A1(add_163_carry_11_), .A2(control_bus[8]), .Z(N113) );
  or02d0 U530 ( .A1(add_163_carry_10_), .A2(n476), .Z(add_163_carry_11_) );
  xn02d1 U531 ( .A1(n476), .A2(add_163_carry_10_), .ZN(N112) );
  or02d0 U532 ( .A1(add_163_carry_9_), .A2(n471), .Z(add_163_carry_10_) );
  xn02d1 U533 ( .A1(n472), .A2(add_163_carry_9_), .ZN(N111) );
  or02d0 U534 ( .A1(add_163_carry_8_), .A2(control_bus[5]), .Z(
        add_163_carry_9_) );
  xn02d1 U535 ( .A1(control_bus[5]), .A2(add_163_carry_8_), .ZN(N110) );
  an02d0 U536 ( .A1(control_bus[4]), .A2(add_163_carry_7_), .Z(
        add_163_carry_8_) );
  xr02d1 U537 ( .A1(add_163_carry_7_), .A2(control_bus[4]), .Z(N109) );
  or02d0 U538 ( .A1(add_163_carry_6_), .A2(control_bus[3]), .Z(
        add_163_carry_7_) );
  xn02d1 U539 ( .A1(control_bus[3]), .A2(add_163_carry_6_), .ZN(N108) );
  or02d0 U540 ( .A1(add_163_carry_5_), .A2(n468), .Z(add_163_carry_6_) );
  xn02d1 U541 ( .A1(n468), .A2(add_163_carry_5_), .ZN(N107) );
  an02d0 U542 ( .A1(N42), .A2(add_163_carry_4_), .Z(add_163_carry_5_) );
  xr02d1 U543 ( .A1(add_163_carry_4_), .A2(N42), .Z(N106) );
  an02d0 U544 ( .A1(n372), .A2(add_163_carry_3_), .Z(add_163_carry_4_) );
  xr02d1 U545 ( .A1(add_163_carry_3_), .A2(n372), .Z(N105) );
  an02d0 U546 ( .A1(n482), .A2(n483), .Z(add_163_carry_3_) );
  xr02d1 U547 ( .A1(n483), .A2(n482), .Z(N104) );
  xr02d1 U548 ( .A1(add_165_carry_15_), .A2(control_bus[12]), .Z(N133) );
  an02d0 U549 ( .A1(control_bus[11]), .A2(add_165_carry_14_), .Z(
        add_165_carry_15_) );
  xr02d1 U550 ( .A1(add_165_carry_14_), .A2(control_bus[11]), .Z(N132) );
  an02d0 U551 ( .A1(n481), .A2(add_165_carry_13_), .Z(add_165_carry_14_) );
  xr02d1 U552 ( .A1(add_165_carry_13_), .A2(n481), .Z(N131) );
  or02d0 U553 ( .A1(add_165_carry_12_), .A2(control_bus[9]), .Z(
        add_165_carry_13_) );
  xn02d1 U554 ( .A1(control_bus[9]), .A2(add_165_carry_12_), .ZN(N130) );
  or02d0 U555 ( .A1(add_165_carry_11_), .A2(control_bus[8]), .Z(
        add_165_carry_12_) );
  xn02d1 U556 ( .A1(control_bus[8]), .A2(add_165_carry_11_), .ZN(N129) );
  or02d0 U557 ( .A1(add_165_carry_10_), .A2(n475), .Z(add_165_carry_11_) );
  xn02d1 U558 ( .A1(n475), .A2(add_165_carry_10_), .ZN(N128) );
  an02d0 U559 ( .A1(n473), .A2(add_165_carry_9_), .Z(add_165_carry_10_) );
  xr02d1 U560 ( .A1(add_165_carry_9_), .A2(n473), .Z(N127) );
  an02d0 U561 ( .A1(control_bus[5]), .A2(add_165_carry_8_), .Z(
        add_165_carry_9_) );
  xr02d1 U562 ( .A1(add_165_carry_8_), .A2(control_bus[5]), .Z(N126) );
  or02d0 U563 ( .A1(add_165_carry_7_), .A2(control_bus[4]), .Z(
        add_165_carry_8_) );
  xn02d1 U564 ( .A1(control_bus[4]), .A2(add_165_carry_7_), .ZN(N125) );
  an02d0 U565 ( .A1(control_bus[3]), .A2(add_165_carry_6_), .Z(
        add_165_carry_7_) );
  xr02d1 U566 ( .A1(add_165_carry_6_), .A2(control_bus[3]), .Z(N124) );
  or02d0 U567 ( .A1(add_165_carry_5_), .A2(n467), .Z(add_165_carry_6_) );
  xn02d1 U568 ( .A1(n467), .A2(add_165_carry_5_), .ZN(N123) );
  or02d0 U569 ( .A1(add_165_carry_4_), .A2(N42), .Z(add_165_carry_5_) );
  xn02d1 U570 ( .A1(N42), .A2(add_165_carry_4_), .ZN(N122) );
  an02d0 U571 ( .A1(n383), .A2(add_165_carry_3_), .Z(add_165_carry_4_) );
  xr02d1 U572 ( .A1(add_165_carry_3_), .A2(n383), .Z(N121) );
  an02d0 U573 ( .A1(n482), .A2(n483), .Z(add_165_carry_3_) );
  xr02d1 U574 ( .A1(n483), .A2(n482), .Z(N120) );
  xr02d1 U575 ( .A1(add_167_carry_15_), .A2(control_bus[12]), .Z(N149) );
  an02d0 U576 ( .A1(control_bus[11]), .A2(add_167_carry_14_), .Z(
        add_167_carry_15_) );
  xr02d1 U577 ( .A1(add_167_carry_14_), .A2(control_bus[11]), .Z(N148) );
  an02d0 U578 ( .A1(n479), .A2(add_167_carry_13_), .Z(add_167_carry_14_) );
  xr02d1 U579 ( .A1(add_167_carry_13_), .A2(n479), .Z(N147) );
  an02d0 U580 ( .A1(control_bus[9]), .A2(add_167_carry_12_), .Z(
        add_167_carry_13_) );
  xr02d1 U581 ( .A1(add_167_carry_12_), .A2(control_bus[9]), .Z(N146) );
  or02d0 U582 ( .A1(add_167_carry_11_), .A2(control_bus[8]), .Z(
        add_167_carry_12_) );
  xn02d1 U583 ( .A1(control_bus[8]), .A2(add_167_carry_11_), .ZN(N145) );
  or02d0 U584 ( .A1(add_167_carry_10_), .A2(n477), .Z(add_167_carry_11_) );
  xn02d1 U585 ( .A1(n477), .A2(add_167_carry_10_), .ZN(N144) );
  an02d0 U586 ( .A1(n473), .A2(add_167_carry_9_), .Z(add_167_carry_10_) );
  xr02d1 U587 ( .A1(add_167_carry_9_), .A2(n473), .Z(N143) );
  an02d0 U588 ( .A1(control_bus[5]), .A2(add_167_carry_8_), .Z(
        add_167_carry_9_) );
  xr02d1 U589 ( .A1(add_167_carry_8_), .A2(control_bus[5]), .Z(N142) );
  an02d0 U590 ( .A1(control_bus[4]), .A2(add_167_carry_7_), .Z(
        add_167_carry_8_) );
  xr02d1 U591 ( .A1(add_167_carry_7_), .A2(control_bus[4]), .Z(N141) );
  an02d0 U592 ( .A1(control_bus[3]), .A2(add_167_carry_6_), .Z(
        add_167_carry_7_) );
  xr02d1 U593 ( .A1(add_167_carry_6_), .A2(control_bus[3]), .Z(N140) );
  or02d0 U594 ( .A1(add_167_carry_5_), .A2(n469), .Z(add_167_carry_6_) );
  xn02d1 U595 ( .A1(n469), .A2(add_167_carry_5_), .ZN(N139) );
  an02d0 U596 ( .A1(N42), .A2(add_167_carry_4_), .Z(add_167_carry_5_) );
  xr02d1 U597 ( .A1(add_167_carry_4_), .A2(N42), .Z(N138) );
  or02d0 U598 ( .A1(add_167_carry_3_), .A2(n363), .Z(add_167_carry_4_) );
  xn02d1 U599 ( .A1(n363), .A2(add_167_carry_3_), .ZN(N137) );
  an02d0 U600 ( .A1(n482), .A2(n483), .Z(add_167_carry_3_) );
  xr02d1 U601 ( .A1(n483), .A2(n482), .Z(N136) );
  xr02d1 U602 ( .A1(add_153_carry_15_), .A2(control_bus[12]), .Z(N37) );
  an02d0 U603 ( .A1(control_bus[11]), .A2(add_153_carry_14_), .Z(
        add_153_carry_15_) );
  xr02d1 U604 ( .A1(add_153_carry_14_), .A2(control_bus[11]), .Z(N36) );
  an02d0 U605 ( .A1(n481), .A2(add_153_carry_13_), .Z(add_153_carry_14_) );
  xr02d1 U606 ( .A1(add_153_carry_13_), .A2(n481), .Z(N35) );
  an02d0 U607 ( .A1(control_bus[9]), .A2(add_153_carry_12_), .Z(
        add_153_carry_13_) );
  xr02d1 U608 ( .A1(add_153_carry_12_), .A2(control_bus[9]), .Z(N34) );
  an02d0 U609 ( .A1(control_bus[8]), .A2(add_153_carry_11_), .Z(
        add_153_carry_12_) );
  xr02d1 U610 ( .A1(add_153_carry_11_), .A2(control_bus[8]), .Z(N33) );
  an02d0 U611 ( .A1(n475), .A2(add_153_carry_10_), .Z(add_153_carry_11_) );
  xr02d1 U612 ( .A1(add_153_carry_10_), .A2(n475), .Z(N32) );
  or02d0 U613 ( .A1(add_153_carry_9_), .A2(n472), .Z(add_153_carry_10_) );
  xn02d1 U614 ( .A1(n472), .A2(add_153_carry_9_), .ZN(N31) );
  or02d0 U615 ( .A1(add_153_carry_8_), .A2(control_bus[5]), .Z(
        add_153_carry_9_) );
  xn02d1 U616 ( .A1(control_bus[5]), .A2(add_153_carry_8_), .ZN(N30) );
  or02d0 U617 ( .A1(add_153_carry_7_), .A2(control_bus[4]), .Z(
        add_153_carry_8_) );
  xn02d1 U618 ( .A1(control_bus[4]), .A2(add_153_carry_7_), .ZN(N29) );
  or02d0 U619 ( .A1(add_153_carry_6_), .A2(control_bus[3]), .Z(
        add_153_carry_7_) );
  xn02d1 U620 ( .A1(control_bus[3]), .A2(add_153_carry_6_), .ZN(N28) );
  an02d0 U621 ( .A1(n467), .A2(add_153_carry_5_), .Z(add_153_carry_6_) );
  xr02d1 U622 ( .A1(add_153_carry_5_), .A2(n467), .Z(N27) );
  or02d0 U623 ( .A1(add_153_carry_4_), .A2(N42), .Z(add_153_carry_5_) );
  xn02d1 U624 ( .A1(N42), .A2(add_153_carry_4_), .ZN(N26) );
  an02d0 U625 ( .A1(n363), .A2(add_153_carry_3_), .Z(add_153_carry_4_) );
  xr02d1 U626 ( .A1(add_153_carry_3_), .A2(n363), .Z(N25) );
  or02d0 U627 ( .A1(n483), .A2(n482), .Z(add_153_carry_3_) );
  xn02d1 U628 ( .A1(n482), .A2(n483), .ZN(N24) );
  inv0d0 U629 ( .I(n483), .ZN(N23) );
  xr02d1 U630 ( .A1(add_155_carry_15_), .A2(control_bus[12]), .Z(N53) );
  or02d0 U631 ( .A1(add_155_carry_14_), .A2(control_bus[11]), .Z(
        add_155_carry_15_) );
  xn02d1 U632 ( .A1(control_bus[11]), .A2(add_155_carry_14_), .ZN(N52) );
  or02d0 U633 ( .A1(add_155_carry_13_), .A2(n479), .Z(add_155_carry_14_) );
  xn02d1 U634 ( .A1(n479), .A2(add_155_carry_13_), .ZN(N51) );
  or02d0 U635 ( .A1(add_155_carry_12_), .A2(control_bus[9]), .Z(
        add_155_carry_13_) );
  xn02d1 U636 ( .A1(control_bus[9]), .A2(add_155_carry_12_), .ZN(N50) );
  or02d0 U637 ( .A1(add_155_carry_11_), .A2(control_bus[8]), .Z(
        add_155_carry_12_) );
  xn02d1 U638 ( .A1(control_bus[8]), .A2(add_155_carry_11_), .ZN(N49) );
  or02d0 U639 ( .A1(add_155_carry_10_), .A2(n477), .Z(add_155_carry_11_) );
  xn02d1 U640 ( .A1(n477), .A2(add_155_carry_10_), .ZN(N48) );
  an02d0 U641 ( .A1(n473), .A2(add_155_carry_9_), .Z(add_155_carry_10_) );
  xr02d1 U642 ( .A1(add_155_carry_9_), .A2(n471), .Z(N47) );
  or02d0 U643 ( .A1(add_155_carry_8_), .A2(control_bus[5]), .Z(
        add_155_carry_9_) );
  xn02d1 U644 ( .A1(control_bus[5]), .A2(add_155_carry_8_), .ZN(N46) );
  an02d0 U645 ( .A1(control_bus[4]), .A2(add_155_carry_7_), .Z(
        add_155_carry_8_) );
  xr02d1 U646 ( .A1(add_155_carry_7_), .A2(control_bus[4]), .Z(N45) );
  or02d0 U647 ( .A1(n467), .A2(control_bus[3]), .Z(add_155_carry_7_) );
  xn02d1 U648 ( .A1(control_bus[3]), .A2(n468), .ZN(N44) );
  inv0d0 U649 ( .I(n468), .ZN(N43) );
  xr02d1 U650 ( .A1(add_157_carry_15_), .A2(control_bus[12]), .Z(N69) );
  an02d0 U651 ( .A1(control_bus[11]), .A2(add_157_carry_14_), .Z(
        add_157_carry_15_) );
  xr02d1 U652 ( .A1(add_157_carry_14_), .A2(control_bus[11]), .Z(N68) );
  or02d0 U653 ( .A1(add_157_carry_13_), .A2(n480), .Z(add_157_carry_14_) );
  xn02d1 U654 ( .A1(n480), .A2(add_157_carry_13_), .ZN(N67) );
  or02d0 U655 ( .A1(add_157_carry_12_), .A2(control_bus[9]), .Z(
        add_157_carry_13_) );
  xn02d1 U656 ( .A1(control_bus[9]), .A2(add_157_carry_12_), .ZN(N66) );
  an02d0 U657 ( .A1(control_bus[8]), .A2(add_157_carry_11_), .Z(
        add_157_carry_12_) );
  xr02d1 U658 ( .A1(add_157_carry_11_), .A2(control_bus[8]), .Z(N65) );
  an02d0 U659 ( .A1(n475), .A2(add_157_carry_10_), .Z(add_157_carry_11_) );
  xr02d1 U660 ( .A1(add_157_carry_10_), .A2(n477), .Z(N64) );
  or02d0 U661 ( .A1(add_157_carry_9_), .A2(n472), .Z(add_157_carry_10_) );
  xn02d1 U662 ( .A1(n472), .A2(add_157_carry_9_), .ZN(N63) );
  or02d0 U663 ( .A1(add_157_carry_8_), .A2(control_bus[5]), .Z(
        add_157_carry_9_) );
  xn02d1 U664 ( .A1(control_bus[5]), .A2(add_157_carry_8_), .ZN(N62) );
  or02d0 U665 ( .A1(add_157_carry_7_), .A2(control_bus[4]), .Z(
        add_157_carry_8_) );
  xn02d1 U666 ( .A1(control_bus[4]), .A2(add_157_carry_7_), .ZN(N61) );
  an02d0 U667 ( .A1(control_bus[3]), .A2(add_157_carry_6_), .Z(
        add_157_carry_7_) );
  xr02d1 U668 ( .A1(add_157_carry_6_), .A2(control_bus[3]), .Z(N60) );
  or02d0 U669 ( .A1(add_157_carry_5_), .A2(n467), .Z(add_157_carry_6_) );
  xn02d1 U670 ( .A1(n469), .A2(add_157_carry_5_), .ZN(N59) );
  or02d0 U671 ( .A1(add_157_carry_4_), .A2(N42), .Z(add_157_carry_5_) );
  xn02d1 U672 ( .A1(N42), .A2(add_157_carry_4_), .ZN(N58) );
  or02d0 U673 ( .A1(n482), .A2(n383), .Z(add_157_carry_4_) );
  xn02d1 U674 ( .A1(n372), .A2(n482), .ZN(N57) );
  inv0d0 U675 ( .I(n482), .ZN(N56) );
  xr02d1 U676 ( .A1(add_159_carry_15_), .A2(control_bus[12]), .Z(N85) );
  an02d0 U677 ( .A1(control_bus[11]), .A2(add_159_carry_14_), .Z(
        add_159_carry_15_) );
  xr02d1 U678 ( .A1(add_159_carry_14_), .A2(control_bus[11]), .Z(N84) );
  an02d0 U679 ( .A1(n479), .A2(add_159_carry_13_), .Z(add_159_carry_14_) );
  xr02d1 U680 ( .A1(add_159_carry_13_), .A2(n479), .Z(N83) );
  or02d0 U681 ( .A1(add_159_carry_12_), .A2(control_bus[9]), .Z(
        add_159_carry_13_) );
  xn02d1 U682 ( .A1(control_bus[9]), .A2(add_159_carry_12_), .ZN(N82) );
  an02d0 U683 ( .A1(control_bus[8]), .A2(add_159_carry_11_), .Z(
        add_159_carry_12_) );
  xr02d1 U684 ( .A1(add_159_carry_11_), .A2(control_bus[8]), .Z(N81) );
  an02d0 U685 ( .A1(n477), .A2(add_159_carry_10_), .Z(add_159_carry_11_) );
  xr02d1 U686 ( .A1(add_159_carry_10_), .A2(n476), .Z(N80) );
  an02d0 U687 ( .A1(n471), .A2(add_159_carry_9_), .Z(add_159_carry_10_) );
  xr02d1 U688 ( .A1(add_159_carry_9_), .A2(n471), .Z(N79) );
  or02d0 U689 ( .A1(add_159_carry_8_), .A2(control_bus[5]), .Z(
        add_159_carry_9_) );
  xn02d1 U690 ( .A1(control_bus[5]), .A2(add_159_carry_8_), .ZN(N78) );
  or02d0 U691 ( .A1(add_159_carry_7_), .A2(control_bus[4]), .Z(
        add_159_carry_8_) );
  xn02d1 U692 ( .A1(control_bus[4]), .A2(add_159_carry_7_), .ZN(N77) );
  or02d0 U693 ( .A1(add_159_carry_6_), .A2(control_bus[3]), .Z(
        add_159_carry_7_) );
  xn02d1 U694 ( .A1(control_bus[3]), .A2(add_159_carry_6_), .ZN(N76) );
  an02d0 U695 ( .A1(n469), .A2(add_159_carry_5_), .Z(add_159_carry_6_) );
  xr02d1 U696 ( .A1(add_159_carry_5_), .A2(n469), .Z(N75) );
  or02d0 U697 ( .A1(add_159_carry_4_), .A2(N42), .Z(add_159_carry_5_) );
  xn02d1 U698 ( .A1(N42), .A2(add_159_carry_4_), .ZN(N74) );
  an02d0 U699 ( .A1(n363), .A2(add_159_carry_3_), .Z(add_159_carry_4_) );
  xr02d1 U700 ( .A1(add_159_carry_3_), .A2(n383), .Z(N73) );
  or02d0 U701 ( .A1(n483), .A2(n482), .Z(add_159_carry_3_) );
  xn02d1 U702 ( .A1(n482), .A2(n483), .ZN(N72) );
  nr03d0 U703 ( .A1(n330), .A2(n327), .A3(n328), .ZN(n364) );
endmodule


module BLENDER_DW_mult_uns_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n742, n744, n746, n748, n749, n750, n751, n755, n756, n758, n759,
         n760, n761, n762, n764, n765, n767, n769, n770, n772, n774, n775,
         n776, n777, n778, n780, n782, n783, n784, n785, n786, n788, n790,
         n791, n792, n793, n794, n796, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n816, n818, n819, n820, n822, n824, n825, n827, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n890, n891, n892, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n956, n957, n958, n959, n960,
         n961, n962, n963, n965, n966, n967;

  nr02d0 U33 ( .A1(n32), .A2(n48), .ZN(product[0]) );
  nr02d0 U34 ( .A1(n49), .A2(n32), .ZN(n65) );
  nr02d0 U35 ( .A1(n50), .A2(n32), .ZN(n66) );
  nr02d0 U36 ( .A1(n51), .A2(n32), .ZN(n67) );
  nr02d0 U37 ( .A1(n52), .A2(n32), .ZN(n68) );
  nr02d0 U38 ( .A1(n53), .A2(n32), .ZN(n69) );
  nr02d0 U39 ( .A1(n54), .A2(n32), .ZN(n70) );
  nr02d0 U40 ( .A1(n55), .A2(n32), .ZN(n71) );
  nr02d0 U41 ( .A1(n56), .A2(n32), .ZN(n72) );
  nr02d0 U42 ( .A1(n57), .A2(n32), .ZN(n73) );
  nr02d0 U43 ( .A1(n58), .A2(n32), .ZN(n74) );
  nr02d0 U44 ( .A1(n59), .A2(n32), .ZN(n75) );
  nr02d0 U45 ( .A1(n60), .A2(n32), .ZN(n76) );
  nr02d0 U46 ( .A1(n61), .A2(n32), .ZN(n77) );
  nr02d0 U47 ( .A1(n62), .A2(n32), .ZN(n78) );
  nr02d0 U48 ( .A1(n63), .A2(n32), .ZN(n79) );
  nr02d0 U49 ( .A1(n33), .A2(n48), .ZN(n80) );
  nr02d0 U50 ( .A1(n33), .A2(n49), .ZN(n81) );
  nr02d0 U51 ( .A1(n50), .A2(n33), .ZN(n82) );
  nr02d0 U52 ( .A1(n51), .A2(n33), .ZN(n83) );
  nr02d0 U53 ( .A1(n52), .A2(n33), .ZN(n84) );
  nr02d0 U54 ( .A1(n53), .A2(n33), .ZN(n85) );
  nr02d0 U55 ( .A1(n54), .A2(n33), .ZN(n86) );
  nr02d0 U56 ( .A1(n55), .A2(n33), .ZN(n87) );
  nr02d0 U57 ( .A1(n56), .A2(n33), .ZN(n88) );
  nr02d0 U58 ( .A1(n57), .A2(n33), .ZN(n89) );
  nr02d0 U59 ( .A1(n58), .A2(n33), .ZN(n90) );
  nr02d0 U60 ( .A1(n59), .A2(n33), .ZN(n91) );
  nr02d0 U61 ( .A1(n60), .A2(n33), .ZN(n92) );
  nr02d0 U62 ( .A1(n61), .A2(n33), .ZN(n93) );
  nr02d0 U63 ( .A1(n62), .A2(n33), .ZN(n94) );
  nr02d0 U64 ( .A1(n63), .A2(n33), .ZN(n95) );
  nr02d0 U65 ( .A1(n34), .A2(n48), .ZN(n96) );
  nr02d0 U66 ( .A1(n34), .A2(n49), .ZN(n97) );
  nr02d0 U67 ( .A1(n34), .A2(n50), .ZN(n98) );
  nr02d0 U68 ( .A1(n51), .A2(n34), .ZN(n99) );
  nr02d0 U69 ( .A1(n52), .A2(n34), .ZN(n100) );
  nr02d0 U70 ( .A1(n53), .A2(n34), .ZN(n101) );
  nr02d0 U71 ( .A1(n54), .A2(n34), .ZN(n102) );
  nr02d0 U72 ( .A1(n55), .A2(n34), .ZN(n103) );
  nr02d0 U73 ( .A1(n56), .A2(n34), .ZN(n104) );
  nr02d0 U74 ( .A1(n57), .A2(n34), .ZN(n105) );
  nr02d0 U75 ( .A1(n58), .A2(n34), .ZN(n106) );
  nr02d0 U76 ( .A1(n59), .A2(n34), .ZN(n107) );
  nr02d0 U77 ( .A1(n60), .A2(n34), .ZN(n108) );
  nr02d0 U78 ( .A1(n61), .A2(n34), .ZN(n109) );
  nr02d0 U79 ( .A1(n62), .A2(n34), .ZN(n110) );
  nr02d0 U80 ( .A1(n63), .A2(n34), .ZN(n111) );
  nr02d0 U81 ( .A1(n35), .A2(n48), .ZN(n112) );
  nr02d0 U82 ( .A1(n35), .A2(n49), .ZN(n113) );
  nr02d0 U83 ( .A1(n35), .A2(n50), .ZN(n114) );
  nr02d0 U84 ( .A1(n35), .A2(n51), .ZN(n115) );
  nr02d0 U85 ( .A1(n52), .A2(n35), .ZN(n116) );
  nr02d0 U86 ( .A1(n53), .A2(n35), .ZN(n117) );
  nr02d0 U87 ( .A1(n54), .A2(n35), .ZN(n118) );
  nr02d0 U88 ( .A1(n55), .A2(n35), .ZN(n119) );
  nr02d0 U89 ( .A1(n56), .A2(n35), .ZN(n120) );
  nr02d0 U90 ( .A1(n57), .A2(n35), .ZN(n121) );
  nr02d0 U91 ( .A1(n58), .A2(n35), .ZN(n122) );
  nr02d0 U92 ( .A1(n59), .A2(n35), .ZN(n123) );
  nr02d0 U93 ( .A1(n60), .A2(n35), .ZN(n124) );
  nr02d0 U94 ( .A1(n61), .A2(n35), .ZN(n125) );
  nr02d0 U95 ( .A1(n62), .A2(n35), .ZN(n126) );
  nr02d0 U96 ( .A1(n63), .A2(n35), .ZN(n127) );
  nr02d0 U97 ( .A1(n36), .A2(n48), .ZN(n128) );
  nr02d0 U98 ( .A1(n36), .A2(n49), .ZN(n129) );
  nr02d0 U99 ( .A1(n36), .A2(n50), .ZN(n130) );
  nr02d0 U100 ( .A1(n36), .A2(n51), .ZN(n131) );
  nr02d0 U101 ( .A1(n36), .A2(n52), .ZN(n132) );
  nr02d0 U102 ( .A1(n53), .A2(n36), .ZN(n133) );
  nr02d0 U103 ( .A1(n54), .A2(n36), .ZN(n134) );
  nr02d0 U104 ( .A1(n55), .A2(n36), .ZN(n135) );
  nr02d0 U105 ( .A1(n56), .A2(n36), .ZN(n136) );
  nr02d0 U106 ( .A1(n57), .A2(n36), .ZN(n137) );
  nr02d0 U107 ( .A1(n58), .A2(n36), .ZN(n138) );
  nr02d0 U108 ( .A1(n59), .A2(n36), .ZN(n139) );
  nr02d0 U109 ( .A1(n60), .A2(n36), .ZN(n140) );
  nr02d0 U110 ( .A1(n61), .A2(n36), .ZN(n141) );
  nr02d0 U111 ( .A1(n62), .A2(n36), .ZN(n142) );
  nr02d0 U112 ( .A1(n63), .A2(n36), .ZN(n143) );
  nr02d0 U113 ( .A1(n37), .A2(n48), .ZN(n144) );
  nr02d0 U114 ( .A1(n37), .A2(n49), .ZN(n145) );
  nr02d0 U115 ( .A1(n37), .A2(n50), .ZN(n146) );
  nr02d0 U116 ( .A1(n37), .A2(n51), .ZN(n147) );
  nr02d0 U117 ( .A1(n37), .A2(n52), .ZN(n148) );
  nr02d0 U118 ( .A1(n37), .A2(n53), .ZN(n149) );
  nr02d0 U119 ( .A1(n54), .A2(n37), .ZN(n150) );
  nr02d0 U120 ( .A1(n55), .A2(n37), .ZN(n151) );
  nr02d0 U121 ( .A1(n37), .A2(n56), .ZN(n152) );
  nr02d0 U122 ( .A1(n57), .A2(n37), .ZN(n153) );
  nr02d0 U123 ( .A1(n58), .A2(n37), .ZN(n154) );
  nr02d0 U124 ( .A1(n59), .A2(n37), .ZN(n155) );
  nr02d0 U125 ( .A1(n60), .A2(n37), .ZN(n156) );
  nr02d0 U126 ( .A1(n61), .A2(n37), .ZN(n157) );
  nr02d0 U127 ( .A1(n62), .A2(n37), .ZN(n158) );
  nr02d0 U128 ( .A1(n63), .A2(n37), .ZN(n159) );
  nr02d0 U129 ( .A1(n38), .A2(n48), .ZN(n160) );
  nr02d0 U130 ( .A1(n38), .A2(n49), .ZN(n161) );
  nr02d0 U131 ( .A1(n38), .A2(n50), .ZN(n162) );
  nr02d0 U132 ( .A1(n38), .A2(n51), .ZN(n163) );
  nr02d0 U133 ( .A1(n38), .A2(n52), .ZN(n164) );
  nr02d0 U134 ( .A1(n38), .A2(n53), .ZN(n165) );
  nr02d0 U135 ( .A1(n38), .A2(n54), .ZN(n166) );
  nr02d0 U136 ( .A1(n55), .A2(n38), .ZN(n167) );
  nr02d0 U137 ( .A1(n38), .A2(n56), .ZN(n168) );
  nr02d0 U138 ( .A1(n57), .A2(n38), .ZN(n169) );
  nr02d0 U139 ( .A1(n58), .A2(n38), .ZN(n170) );
  nr02d0 U140 ( .A1(n59), .A2(n38), .ZN(n171) );
  nr02d0 U141 ( .A1(n60), .A2(n38), .ZN(n172) );
  nr02d0 U142 ( .A1(n61), .A2(n38), .ZN(n173) );
  nr02d0 U143 ( .A1(n62), .A2(n38), .ZN(n174) );
  nr02d0 U144 ( .A1(n63), .A2(n38), .ZN(n175) );
  nr02d0 U145 ( .A1(n39), .A2(n48), .ZN(n176) );
  nr02d0 U146 ( .A1(n39), .A2(n49), .ZN(n177) );
  nr02d0 U147 ( .A1(n39), .A2(n50), .ZN(n178) );
  nr02d0 U148 ( .A1(n39), .A2(n51), .ZN(n179) );
  nr02d0 U149 ( .A1(n39), .A2(n52), .ZN(n180) );
  nr02d0 U150 ( .A1(n39), .A2(n53), .ZN(n181) );
  nr02d0 U151 ( .A1(n39), .A2(n54), .ZN(n182) );
  nr02d0 U152 ( .A1(n39), .A2(n55), .ZN(n183) );
  nr02d0 U153 ( .A1(n39), .A2(n56), .ZN(n184) );
  nr02d0 U154 ( .A1(n39), .A2(n57), .ZN(n185) );
  nr02d0 U155 ( .A1(n58), .A2(n39), .ZN(n186) );
  nr02d0 U156 ( .A1(n59), .A2(n39), .ZN(n187) );
  nr02d0 U157 ( .A1(n60), .A2(n39), .ZN(n188) );
  nr02d0 U158 ( .A1(n61), .A2(n39), .ZN(n189) );
  nr02d0 U159 ( .A1(n62), .A2(n39), .ZN(n190) );
  nr02d0 U160 ( .A1(n63), .A2(n39), .ZN(n191) );
  nr02d0 U161 ( .A1(n40), .A2(n48), .ZN(n192) );
  nr02d0 U162 ( .A1(n40), .A2(n49), .ZN(n193) );
  nr02d0 U163 ( .A1(n40), .A2(n50), .ZN(n194) );
  nr02d0 U164 ( .A1(n40), .A2(n51), .ZN(n195) );
  nr02d0 U165 ( .A1(n40), .A2(n52), .ZN(n196) );
  nr02d0 U166 ( .A1(n53), .A2(n40), .ZN(n197) );
  nr02d0 U167 ( .A1(n54), .A2(n40), .ZN(n198) );
  nr02d0 U168 ( .A1(n55), .A2(n40), .ZN(n199) );
  nr02d0 U169 ( .A1(n56), .A2(n40), .ZN(n200) );
  nr02d0 U170 ( .A1(n57), .A2(n40), .ZN(n201) );
  nr02d0 U171 ( .A1(n58), .A2(n40), .ZN(n202) );
  nr02d0 U172 ( .A1(n59), .A2(n40), .ZN(n203) );
  nr02d0 U173 ( .A1(n60), .A2(n40), .ZN(n204) );
  nr02d0 U174 ( .A1(n61), .A2(n40), .ZN(n205) );
  nr02d0 U175 ( .A1(n62), .A2(n40), .ZN(n206) );
  nr02d0 U176 ( .A1(n63), .A2(n40), .ZN(n207) );
  nr02d0 U177 ( .A1(n41), .A2(n48), .ZN(n208) );
  nr02d0 U178 ( .A1(n41), .A2(n49), .ZN(n209) );
  nr02d0 U179 ( .A1(n41), .A2(n50), .ZN(n210) );
  nr02d0 U180 ( .A1(n41), .A2(n51), .ZN(n211) );
  nr02d0 U181 ( .A1(n41), .A2(n52), .ZN(n212) );
  nr02d0 U182 ( .A1(n41), .A2(n53), .ZN(n213) );
  nr02d0 U183 ( .A1(n41), .A2(n54), .ZN(n214) );
  nr02d0 U184 ( .A1(n55), .A2(n41), .ZN(n215) );
  nr02d0 U185 ( .A1(n41), .A2(n56), .ZN(n216) );
  nr02d0 U186 ( .A1(n57), .A2(n41), .ZN(n217) );
  nr02d0 U187 ( .A1(n58), .A2(n41), .ZN(n218) );
  nr02d0 U188 ( .A1(n59), .A2(n41), .ZN(n219) );
  nr02d0 U189 ( .A1(n60), .A2(n41), .ZN(n220) );
  nr02d0 U190 ( .A1(n61), .A2(n41), .ZN(n221) );
  nr02d0 U191 ( .A1(n62), .A2(n41), .ZN(n222) );
  nr02d0 U192 ( .A1(n63), .A2(n41), .ZN(n223) );
  nr02d0 U193 ( .A1(n42), .A2(n48), .ZN(n224) );
  nr02d0 U194 ( .A1(n42), .A2(n49), .ZN(n225) );
  nr02d0 U195 ( .A1(n42), .A2(n50), .ZN(n226) );
  nr02d0 U196 ( .A1(n42), .A2(n51), .ZN(n227) );
  nr02d0 U197 ( .A1(n42), .A2(n52), .ZN(n228) );
  nr02d0 U198 ( .A1(n42), .A2(n53), .ZN(n229) );
  nr02d0 U199 ( .A1(n42), .A2(n54), .ZN(n230) );
  nr02d0 U200 ( .A1(n42), .A2(n55), .ZN(n231) );
  nr02d0 U201 ( .A1(n42), .A2(n56), .ZN(n232) );
  nr02d0 U202 ( .A1(n42), .A2(n57), .ZN(n233) );
  nr02d0 U203 ( .A1(n42), .A2(n58), .ZN(n234) );
  nr02d0 U204 ( .A1(n59), .A2(n42), .ZN(n235) );
  nr02d0 U205 ( .A1(n60), .A2(n42), .ZN(n236) );
  nr02d0 U206 ( .A1(n61), .A2(n42), .ZN(n237) );
  nr02d0 U207 ( .A1(n62), .A2(n42), .ZN(n238) );
  nr02d0 U208 ( .A1(n63), .A2(n42), .ZN(n239) );
  nr02d0 U209 ( .A1(n43), .A2(n48), .ZN(n240) );
  nr02d0 U210 ( .A1(n43), .A2(n49), .ZN(n241) );
  nr02d0 U211 ( .A1(n43), .A2(n50), .ZN(n242) );
  nr02d0 U212 ( .A1(n43), .A2(n51), .ZN(n243) );
  nr02d0 U213 ( .A1(n43), .A2(n52), .ZN(n244) );
  nr02d0 U214 ( .A1(n43), .A2(n53), .ZN(n245) );
  nr02d0 U215 ( .A1(n43), .A2(n54), .ZN(n246) );
  nr02d0 U216 ( .A1(n43), .A2(n55), .ZN(n247) );
  nr02d0 U217 ( .A1(n43), .A2(n56), .ZN(n248) );
  nr02d0 U218 ( .A1(n43), .A2(n57), .ZN(n249) );
  nr02d0 U219 ( .A1(n43), .A2(n58), .ZN(n250) );
  nr02d0 U220 ( .A1(n59), .A2(n43), .ZN(n251) );
  nr02d0 U221 ( .A1(n60), .A2(n43), .ZN(n252) );
  nr02d0 U222 ( .A1(n61), .A2(n43), .ZN(n253) );
  nr02d0 U223 ( .A1(n62), .A2(n43), .ZN(n254) );
  nr02d0 U224 ( .A1(n63), .A2(n43), .ZN(n255) );
  nr02d0 U225 ( .A1(n44), .A2(n48), .ZN(n256) );
  nr02d0 U226 ( .A1(n44), .A2(n49), .ZN(n257) );
  nr02d0 U227 ( .A1(n44), .A2(n50), .ZN(n258) );
  nr02d0 U228 ( .A1(n44), .A2(n51), .ZN(n259) );
  nr02d0 U229 ( .A1(n44), .A2(n52), .ZN(n260) );
  nr02d0 U230 ( .A1(n44), .A2(n53), .ZN(n261) );
  nr02d0 U231 ( .A1(n44), .A2(n54), .ZN(n262) );
  nr02d0 U232 ( .A1(n44), .A2(n55), .ZN(n263) );
  nr02d0 U233 ( .A1(n44), .A2(n56), .ZN(n264) );
  nr02d0 U234 ( .A1(n44), .A2(n57), .ZN(n265) );
  nr02d0 U235 ( .A1(n44), .A2(n58), .ZN(n266) );
  nr02d0 U236 ( .A1(n44), .A2(n59), .ZN(n267) );
  nr02d0 U237 ( .A1(n60), .A2(n44), .ZN(n268) );
  nr02d0 U238 ( .A1(n61), .A2(n44), .ZN(n269) );
  nr02d0 U239 ( .A1(n62), .A2(n44), .ZN(n270) );
  nr02d0 U240 ( .A1(n63), .A2(n44), .ZN(n271) );
  nr02d0 U241 ( .A1(n45), .A2(n48), .ZN(n272) );
  nr02d0 U242 ( .A1(n45), .A2(n49), .ZN(n273) );
  nr02d0 U243 ( .A1(n45), .A2(n50), .ZN(n274) );
  nr02d0 U244 ( .A1(n45), .A2(n51), .ZN(n275) );
  nr02d0 U245 ( .A1(n45), .A2(n52), .ZN(n276) );
  nr02d0 U246 ( .A1(n45), .A2(n53), .ZN(n277) );
  nr02d0 U247 ( .A1(n45), .A2(n54), .ZN(n278) );
  nr02d0 U248 ( .A1(n45), .A2(n55), .ZN(n279) );
  nr02d0 U249 ( .A1(n45), .A2(n56), .ZN(n280) );
  nr02d0 U250 ( .A1(n45), .A2(n57), .ZN(n281) );
  nr02d0 U251 ( .A1(n45), .A2(n58), .ZN(n282) );
  nr02d0 U252 ( .A1(n45), .A2(n59), .ZN(n283) );
  nr02d0 U253 ( .A1(n45), .A2(n60), .ZN(n284) );
  nr02d0 U254 ( .A1(n61), .A2(n45), .ZN(n285) );
  nr02d0 U255 ( .A1(n62), .A2(n45), .ZN(n286) );
  nr02d0 U256 ( .A1(n63), .A2(n45), .ZN(n287) );
  nr02d0 U257 ( .A1(n46), .A2(n48), .ZN(n288) );
  nr02d0 U258 ( .A1(n46), .A2(n49), .ZN(n289) );
  nr02d0 U259 ( .A1(n46), .A2(n50), .ZN(n290) );
  nr02d0 U260 ( .A1(n46), .A2(n51), .ZN(n291) );
  nr02d0 U261 ( .A1(n46), .A2(n52), .ZN(n292) );
  nr02d0 U262 ( .A1(n46), .A2(n53), .ZN(n293) );
  nr02d0 U263 ( .A1(n46), .A2(n54), .ZN(n294) );
  nr02d0 U264 ( .A1(n46), .A2(n55), .ZN(n295) );
  nr02d0 U265 ( .A1(n46), .A2(n56), .ZN(n296) );
  nr02d0 U266 ( .A1(n46), .A2(n57), .ZN(n297) );
  nr02d0 U267 ( .A1(n46), .A2(n58), .ZN(n298) );
  nr02d0 U268 ( .A1(n46), .A2(n59), .ZN(n299) );
  nr02d0 U269 ( .A1(n46), .A2(n60), .ZN(n300) );
  nr02d0 U270 ( .A1(n46), .A2(n61), .ZN(n301) );
  nr02d0 U271 ( .A1(n62), .A2(n46), .ZN(n302) );
  nr02d0 U272 ( .A1(n63), .A2(n46), .ZN(n303) );
  nr02d0 U273 ( .A1(n47), .A2(n48), .ZN(n304) );
  nr02d0 U274 ( .A1(n47), .A2(n49), .ZN(n305) );
  nr02d0 U275 ( .A1(n47), .A2(n50), .ZN(n306) );
  nr02d0 U276 ( .A1(n47), .A2(n51), .ZN(n307) );
  nr02d0 U277 ( .A1(n47), .A2(n52), .ZN(n308) );
  nr02d0 U278 ( .A1(n47), .A2(n53), .ZN(n309) );
  nr02d0 U279 ( .A1(n47), .A2(n54), .ZN(n310) );
  nr02d0 U280 ( .A1(n47), .A2(n55), .ZN(n311) );
  nr02d0 U281 ( .A1(n47), .A2(n56), .ZN(n312) );
  nr02d0 U282 ( .A1(n47), .A2(n57), .ZN(n313) );
  nr02d0 U283 ( .A1(n47), .A2(n58), .ZN(n314) );
  nr02d0 U284 ( .A1(n47), .A2(n59), .ZN(n315) );
  nr02d0 U285 ( .A1(n47), .A2(n60), .ZN(n316) );
  nr02d0 U286 ( .A1(n47), .A2(n61), .ZN(n317) );
  nr02d0 U287 ( .A1(n62), .A2(n47), .ZN(n318) );
  nr02d0 U288 ( .A1(n63), .A2(n47), .ZN(n319) );
  ah01d0 U289 ( .A(n81), .B(n66), .CO(n321), .S(n320) );
  ah01d0 U290 ( .A(n82), .B(n97), .CO(n323), .S(n322) );
  ah01d0 U292 ( .A(n98), .B(n83), .CO(n327), .S(n326) );
  ah01d0 U295 ( .A(n99), .B(n114), .CO(n333), .S(n332) );
  ah01d0 U299 ( .A(n115), .B(n100), .CO(n341), .S(n340) );
  ah01d0 U304 ( .A(n116), .B(n131), .CO(n351), .S(n350) );
  ah01d0 U310 ( .A(n132), .B(n351), .CO(n363), .S(n362) );
  ah01d0 U317 ( .A(n193), .B(n88), .CO(n377), .S(n376) );
  ah01d0 U325 ( .A(n194), .B(n104), .CO(n393), .S(n392) );
  ah01d0 U334 ( .A(n195), .B(n120), .CO(n411), .S(n410) );
  ah01d0 U344 ( .A(n196), .B(n136), .CO(n431), .S(n430) );
  ah01d0 U355 ( .A(n197), .B(n152), .CO(n453), .S(n452) );
  ah01d0 U367 ( .A(n198), .B(n168), .CO(n477), .S(n476) );
  ah01d0 U380 ( .A(n214), .B(n169), .CO(n503), .S(n502) );
  ah01d0 U394 ( .A(n200), .B(n215), .CO(n531), .S(n530) );
  nd02d1 U499 ( .A1(n80), .A2(n65), .ZN(n767) );
  nd02d1 U505 ( .A1(n320), .A2(n96), .ZN(n770) );
  nd02d1 U508 ( .A1(n960), .A2(n770), .ZN(n895) );
  xn02d1 U512 ( .A1(n895), .A2(n769), .ZN(product[2]) );
  nd02d1 U513 ( .A1(n324), .A2(n322), .ZN(n775) );
  nr02d0 U514 ( .A1(n324), .A2(n322), .ZN(n776) );
  nd02d1 U516 ( .A1(n742), .A2(n775), .ZN(n896) );
  oai21d1 U517 ( .B1(n776), .B2(n774), .A(n775), .ZN(n777) );
  xr02d1 U518 ( .A1(n896), .A2(n774), .Z(product[3]) );
  nd02d1 U519 ( .A1(n330), .A2(n328), .ZN(n778) );
  nd02d1 U522 ( .A1(n962), .A2(n778), .ZN(n897) );
  xn02d1 U526 ( .A1(n897), .A2(n777), .ZN(product[4]) );
  nd02d1 U527 ( .A1(n338), .A2(n336), .ZN(n783) );
  nr02d0 U528 ( .A1(n338), .A2(n336), .ZN(n784) );
  nd02d1 U530 ( .A1(n744), .A2(n783), .ZN(n898) );
  oai21d1 U531 ( .B1(n784), .B2(n782), .A(n783), .ZN(n785) );
  xr02d1 U532 ( .A1(n898), .A2(n782), .Z(product[5]) );
  nd02d1 U533 ( .A1(n348), .A2(n346), .ZN(n786) );
  nd02d1 U536 ( .A1(n961), .A2(n786), .ZN(n899) );
  xn02d1 U540 ( .A1(n899), .A2(n785), .ZN(product[6]) );
  nd02d1 U541 ( .A1(n360), .A2(n358), .ZN(n791) );
  nr02d0 U542 ( .A1(n360), .A2(n358), .ZN(n792) );
  nd02d1 U544 ( .A1(n746), .A2(n791), .ZN(n900) );
  oai21d1 U545 ( .B1(n792), .B2(n790), .A(n791), .ZN(n793) );
  xr02d1 U546 ( .A1(n900), .A2(n790), .Z(product[7]) );
  nd02d1 U547 ( .A1(n374), .A2(n361), .ZN(n794) );
  nd02d1 U550 ( .A1(n959), .A2(n794), .ZN(n901) );
  xn02d1 U554 ( .A1(n901), .A2(n793), .ZN(product[8]) );
  nd02d1 U555 ( .A1(n390), .A2(n375), .ZN(n799) );
  nr02d0 U556 ( .A1(n390), .A2(n375), .ZN(n800) );
  nd02d1 U558 ( .A1(n748), .A2(n799), .ZN(n902) );
  oai21d1 U559 ( .B1(n798), .B2(n800), .A(n799), .ZN(n801) );
  xr02d1 U561 ( .A1(n798), .A2(n902), .Z(product[9]) );
  nd02d1 U562 ( .A1(n408), .A2(n391), .ZN(n803) );
  nr02d0 U563 ( .A1(n408), .A2(n391), .ZN(n804) );
  nd02d1 U565 ( .A1(n749), .A2(n803), .ZN(n903) );
  oai21d1 U566 ( .B1(n802), .B2(n804), .A(n803), .ZN(n805) );
  xr02d1 U567 ( .A1(n802), .A2(n903), .Z(product[10]) );
  nd02d1 U568 ( .A1(n428), .A2(n409), .ZN(n806) );
  nr02d0 U569 ( .A1(n428), .A2(n409), .ZN(n807) );
  nd02d1 U571 ( .A1(n750), .A2(n806), .ZN(n904) );
  oai21d1 U572 ( .B1(n807), .B2(n803), .A(n806), .ZN(n808) );
  nr02d0 U573 ( .A1(n807), .A2(n804), .ZN(n809) );
  xn02d1 U575 ( .A1(n805), .A2(n904), .ZN(product[11]) );
  nd02d1 U576 ( .A1(n450), .A2(n429), .ZN(n811) );
  nr02d0 U577 ( .A1(n450), .A2(n429), .ZN(n812) );
  nd02d1 U579 ( .A1(n751), .A2(n811), .ZN(n905) );
  oai21d1 U580 ( .B1(n810), .B2(n812), .A(n811), .ZN(n813) );
  xr02d1 U581 ( .A1(n810), .A2(n905), .Z(product[12]) );
  nd02d1 U582 ( .A1(n474), .A2(n451), .ZN(n814) );
  nd02d1 U585 ( .A1(n958), .A2(n814), .ZN(n906) );
  xn02d1 U590 ( .A1(n813), .A2(n906), .ZN(product[13]) );
  nd02d1 U591 ( .A1(n500), .A2(n475), .ZN(n820) );
  nd02d1 U594 ( .A1(n956), .A2(n820), .ZN(n907) );
  xn02d1 U598 ( .A1(n819), .A2(n907), .ZN(product[14]) );
  nd02d1 U599 ( .A1(n528), .A2(n501), .ZN(n825) );
  nd02d1 U602 ( .A1(n957), .A2(n825), .ZN(n908) );
  nd02d1 U606 ( .A1(n957), .A2(n956), .ZN(n830) );
  oai21d1 U607 ( .B1(n830), .B2(n818), .A(n829), .ZN(n831) );
  xr02d1 U609 ( .A1(n824), .A2(n908), .Z(product[15]) );
  nd02d1 U610 ( .A1(n556), .A2(n529), .ZN(n833) );
  nr02d0 U611 ( .A1(n556), .A2(n529), .ZN(n834) );
  nd02d1 U613 ( .A1(n755), .A2(n833), .ZN(n909) );
  oai21d1 U614 ( .B1(n832), .B2(n834), .A(n833), .ZN(n835) );
  xr02d1 U615 ( .A1(n832), .A2(n909), .Z(product[16]) );
  nd02d1 U616 ( .A1(n582), .A2(n557), .ZN(n836) );
  nr02d0 U617 ( .A1(n582), .A2(n557), .ZN(n837) );
  nd02d1 U619 ( .A1(n756), .A2(n836), .ZN(n910) );
  oai21d1 U620 ( .B1(n837), .B2(n833), .A(n836), .ZN(n838) );
  nr02d0 U621 ( .A1(n837), .A2(n834), .ZN(n839) );
  xn02d1 U624 ( .A1(n835), .A2(n910), .ZN(product[17]) );
  nd02d1 U625 ( .A1(n606), .A2(n583), .ZN(n842) );
  nr02d0 U626 ( .A1(n606), .A2(n583), .ZN(n843) );
  nd02d1 U628 ( .A1(n845), .A2(n842), .ZN(n911) );
  xn02d1 U632 ( .A1(n841), .A2(n911), .ZN(product[18]) );
  nd02d1 U633 ( .A1(n628), .A2(n607), .ZN(n847) );
  nr02d0 U634 ( .A1(n628), .A2(n607), .ZN(n848) );
  nd02d1 U636 ( .A1(n758), .A2(n847), .ZN(n912) );
  oai21d1 U637 ( .B1(n848), .B2(n842), .A(n847), .ZN(n849) );
  nr02d0 U638 ( .A1(n848), .A2(n843), .ZN(n850) );
  nd02d1 U641 ( .A1(n648), .A2(n629), .ZN(n852) );
  nr02d0 U642 ( .A1(n648), .A2(n629), .ZN(n853) );
  nd02d1 U644 ( .A1(n759), .A2(n852), .ZN(n913) );
  oai21d1 U645 ( .B1(n851), .B2(n853), .A(n852), .ZN(n854) );
  xr02d1 U646 ( .A1(n851), .A2(n913), .Z(product[20]) );
  nd02d1 U647 ( .A1(n666), .A2(n649), .ZN(n855) );
  nr02d0 U648 ( .A1(n666), .A2(n649), .ZN(n856) );
  nd02d1 U650 ( .A1(n760), .A2(n855), .ZN(n914) );
  oai21d1 U651 ( .B1(n856), .B2(n852), .A(n855), .ZN(n857) );
  nr02d0 U652 ( .A1(n853), .A2(n856), .ZN(n858) );
  nd02d1 U654 ( .A1(n850), .A2(n858), .ZN(n860) );
  oai21d1 U655 ( .B1(n840), .B2(n860), .A(n859), .ZN(n861) );
  xn02d1 U657 ( .A1(n854), .A2(n914), .ZN(product[21]) );
  nd02d1 U658 ( .A1(n682), .A2(n667), .ZN(n863) );
  nr02d0 U659 ( .A1(n682), .A2(n667), .ZN(n864) );
  nd02d1 U661 ( .A1(n761), .A2(n863), .ZN(n915) );
  oai21d1 U662 ( .B1(n862), .B2(n864), .A(n863), .ZN(n865) );
  xr02d1 U663 ( .A1(n862), .A2(n915), .Z(product[22]) );
  nd02d1 U664 ( .A1(n696), .A2(n683), .ZN(n866) );
  nr02d0 U665 ( .A1(n696), .A2(n683), .ZN(n867) );
  nd02d1 U667 ( .A1(n762), .A2(n866), .ZN(n916) );
  oai21d1 U668 ( .B1(n867), .B2(n863), .A(n866), .ZN(n868) );
  nr02d0 U669 ( .A1(n864), .A2(n867), .ZN(n869) );
  oai21d1 U672 ( .B1(n862), .B2(n871), .A(n870), .ZN(n872) );
  xn02d1 U673 ( .A1(n865), .A2(n916), .ZN(product[23]) );
  nd02d1 U674 ( .A1(n708), .A2(n697), .ZN(n873) );
  nr02d0 U675 ( .A1(n708), .A2(n697), .ZN(n874) );
  nd02d1 U677 ( .A1(n876), .A2(n873), .ZN(n917) );
  xn02d1 U681 ( .A1(n872), .A2(n917), .ZN(product[24]) );
  nd02d1 U682 ( .A1(n718), .A2(n709), .ZN(n878) );
  nr02d0 U683 ( .A1(n718), .A2(n709), .ZN(n879) );
  nd02d1 U685 ( .A1(n764), .A2(n878), .ZN(n918) );
  oai21d1 U686 ( .B1(n873), .B2(n879), .A(n878), .ZN(n880) );
  nr02d0 U687 ( .A1(n874), .A2(n879), .ZN(n881) );
  nd02d1 U689 ( .A1(n869), .A2(n881), .ZN(n883) );
  oai21d1 U690 ( .B1(n862), .B2(n883), .A(n882), .ZN(n884) );
  nd02d1 U692 ( .A1(n726), .A2(n719), .ZN(n885) );
  nr02d0 U693 ( .A1(n726), .A2(n719), .ZN(n886) );
  nd02d1 U695 ( .A1(n765), .A2(n885), .ZN(n919) );
  oai21d1 U696 ( .B1(n882), .B2(n886), .A(n885), .ZN(n887) );
  nr02d0 U697 ( .A1(n883), .A2(n886), .ZN(n888) );
  xn02d1 U699 ( .A1(n884), .A2(n919), .ZN(product[26]) );
  ad01d0 U708 ( .A(n727), .B(n732), .CI(n967), .CO(n890), .S(product[27]) );
  or02d1 U709 ( .A1(n500), .A2(n475), .Z(n956) );
  or02d1 U710 ( .A1(n528), .A2(n501), .Z(n957) );
  or02d1 U711 ( .A1(n474), .A2(n451), .Z(n958) );
  or02d1 U712 ( .A1(n374), .A2(n361), .Z(n959) );
  or02d1 U713 ( .A1(n320), .A2(n96), .Z(n960) );
  or02d1 U714 ( .A1(n348), .A2(n346), .Z(n961) );
  or02d1 U715 ( .A1(n330), .A2(n328), .Z(n962) );
  or02d1 U716 ( .A1(n80), .A2(n65), .Z(n963) );
  an02d1 U717 ( .A1(n963), .A2(n767), .Z(product[1]) );
  aoi21d1 U718 ( .B1(n809), .B2(n801), .A(n808), .ZN(n810) );
  xn02d1 U719 ( .A1(n965), .A2(n912), .ZN(product[19]) );
  aor21d1 U720 ( .B1(n841), .B2(n845), .A(n844), .Z(n965) );
  xn02d1 U721 ( .A1(n966), .A2(n918), .ZN(product[25]) );
  aor21d1 U722 ( .B1(n872), .B2(n876), .A(n875), .Z(n966) );
  ad01d0 U723 ( .A(n416), .B(n403), .CI(n418), .CO(n425), .S(n424) );
  ad01d0 U724 ( .A(n345), .B(n352), .CI(n354), .CO(n359), .S(n358) );
  ad01d0 U725 ( .A(n423), .B(n438), .CI(n440), .CO(n447), .S(n446) );
  ad01d0 U726 ( .A(n385), .B(n396), .CI(n398), .CO(n405), .S(n404) );
  ad01d0 U727 ( .A(n413), .B(n415), .CI(n417), .CO(n439), .S(n438) );
  ad01d0 U728 ( .A(n503), .B(n530), .CI(n505), .CO(n535), .S(n534) );
  ad01d0 U729 ( .A(n359), .B(n370), .CI(n372), .CO(n375), .S(n374) );
  ad01d0 U730 ( .A(n473), .B(n496), .CI(n498), .CO(n501), .S(n500) );
  ad01d0 U731 ( .A(n407), .B(n424), .CI(n426), .CO(n429), .S(n428) );
  ad01d0 U732 ( .A(n449), .B(n470), .CI(n472), .CO(n475), .S(n474) );
  ad01d0 U733 ( .A(n427), .B(n446), .CI(n448), .CO(n451), .S(n450) );
  ad01d0 U734 ( .A(n555), .B(n578), .CI(n580), .CO(n583), .S(n582) );
  ad01d0 U735 ( .A(n692), .B(n681), .CI(n694), .CO(n697), .S(n696) );
  ad01d0 U736 ( .A(n389), .B(n404), .CI(n406), .CO(n409), .S(n408) );
  ad01d0 U737 ( .A(n527), .B(n552), .CI(n554), .CO(n557), .S(n556) );
  ad01d0 U738 ( .A(n602), .B(n581), .CI(n604), .CO(n607), .S(n606) );
  ad01d0 U739 ( .A(n644), .B(n627), .CI(n646), .CO(n649), .S(n648) );
  ad01d0 U740 ( .A(n678), .B(n665), .CI(n680), .CO(n683), .S(n682) );
  ad01d0 U741 ( .A(n704), .B(n695), .CI(n706), .CO(n709), .S(n708) );
  ad01d0 U742 ( .A(n373), .B(n386), .CI(n388), .CO(n391), .S(n390) );
  ad01d0 U743 ( .A(n499), .B(n524), .CI(n526), .CO(n529), .S(n528) );
  ad01d0 U744 ( .A(n624), .B(n605), .CI(n626), .CO(n629), .S(n628) );
  ad01d0 U745 ( .A(n662), .B(n647), .CI(n664), .CO(n667), .S(n666) );
  ad01d0 U746 ( .A(n382), .B(n371), .CI(n384), .CO(n389), .S(n388) );
  ad01d0 U747 ( .A(n577), .B(n600), .CI(n579), .CO(n605), .S(n604) );
  ad01d0 U748 ( .A(n623), .B(n642), .CI(n625), .CO(n647), .S(n646) );
  ad01d0 U749 ( .A(n601), .B(n622), .CI(n603), .CO(n627), .S(n626) );
  ad01d0 U750 ( .A(n454), .B(n437), .CI(n456), .CO(n463), .S(n462) );
  aor21d1 U751 ( .B1(n861), .B2(n888), .A(n887), .Z(n967) );
  ad01d0 U752 ( .A(n736), .B(n733), .CI(n890), .CO(n891), .S(product[28]) );
  ad01d0 U753 ( .A(n284), .B(n269), .CI(n299), .CO(n711), .S(n710) );
  ad01d0 U754 ( .A(n145), .B(n70), .CI(n340), .CO(n345), .S(n344) );
  ad01d0 U755 ( .A(n341), .B(n101), .CI(n146), .CO(n353), .S(n352) );
  ad01d0 U756 ( .A(n243), .B(n123), .CI(n478), .CO(n485), .S(n484) );
  ad01d0 U757 ( .A(n165), .B(n150), .CI(n393), .CO(n413), .S(n412) );
  ad01d0 U758 ( .A(n479), .B(n244), .CI(n481), .CO(n509), .S(n508) );
  ad01d0 U759 ( .A(n154), .B(n229), .CI(n502), .CO(n507), .S(n506) );
  ad01d0 U760 ( .A(n245), .B(n155), .CI(n507), .CO(n537), .S(n536) );
  ad01d0 U761 ( .A(n631), .B(n220), .CI(n280), .CO(n653), .S(n652) );
  ad01d0 U762 ( .A(n630), .B(n279), .CI(n611), .CO(n635), .S(n634) );
  ad01d0 U763 ( .A(n172), .B(n563), .CI(n586), .CO(n591), .S(n590) );
  ad01d0 U764 ( .A(n281), .B(n651), .CI(n221), .CO(n671), .S(n670) );
  ad01d0 U765 ( .A(n353), .B(n355), .CI(n364), .CO(n371), .S(n370) );
  ad01d0 U766 ( .A(n516), .B(n495), .CI(n518), .CO(n525), .S(n524) );
  ad01d0 U767 ( .A(n595), .B(n597), .CI(n616), .CO(n623), .S(n622) );
  ad01d0 U768 ( .A(n571), .B(n573), .CI(n594), .CO(n601), .S(n600) );
  ad01d0 U769 ( .A(n617), .B(n636), .CI(n619), .CO(n643), .S(n642) );
  ad01d0 U770 ( .A(n489), .B(n512), .CI(n289), .CO(n519), .S(n518) );
  ad01d0 U771 ( .A(n430), .B(n106), .CI(n226), .CO(n437), .S(n436) );
  ad01d0 U772 ( .A(n210), .B(n105), .CI(n180), .CO(n415), .S(n414) );
  ad01d0 U773 ( .A(n431), .B(n212), .CI(n182), .CO(n455), .S(n454) );
  ad01d0 U774 ( .A(n185), .B(n170), .CI(n230), .CO(n533), .S(n532) );
  ad01d0 U775 ( .A(n535), .B(n261), .CI(n156), .CO(n565), .S(n564) );
  ad01d0 U776 ( .A(n267), .B(n252), .CI(n282), .CO(n685), .S(n684) );
  ad01d0 U777 ( .A(n130), .B(n333), .CI(n85), .CO(n343), .S(n342) );
  ad01d0 U778 ( .A(n217), .B(n202), .CI(n232), .CO(n585), .S(n584) );
  ad01d0 U779 ( .A(n668), .B(n296), .CI(n653), .CO(n673), .S(n672) );
  ad01d0 U780 ( .A(n234), .B(n249), .CI(n219), .CO(n631), .S(n630) );
  ad01d0 U781 ( .A(n584), .B(n262), .CI(n561), .CO(n589), .S(n588) );
  ad01d0 U782 ( .A(n251), .B(n266), .CI(n236), .CO(n669), .S(n668) );
  ad01d0 U783 ( .A(n669), .B(n237), .CI(n297), .CO(n687), .S(n686) );
  ad01d0 U784 ( .A(n485), .B(n508), .CI(n274), .CO(n515), .S(n514) );
  ad01d0 U785 ( .A(n86), .B(n161), .CI(n350), .CO(n355), .S(n354) );
  ad01d0 U786 ( .A(n241), .B(n432), .CI(n434), .CO(n441), .S(n440) );
  ad01d0 U787 ( .A(n378), .B(n369), .CI(n380), .CO(n387), .S(n386) );
  ad01d0 U788 ( .A(n465), .B(n93), .CI(n486), .CO(n493), .S(n492) );
  ad01d0 U789 ( .A(n171), .B(n533), .CI(n558), .CO(n563), .S(n562) );
  ad01d0 U790 ( .A(n587), .B(n188), .CI(n608), .CO(n613), .S(n612) );
  ad01d0 U791 ( .A(n487), .B(n109), .CI(n510), .CO(n517), .S(n516) );
  ad01d0 U792 ( .A(n544), .B(n523), .CI(n546), .CO(n553), .S(n552) );
  ad01d0 U793 ( .A(n90), .B(n225), .CI(n397), .CO(n419), .S(n418) );
  ad01d0 U794 ( .A(n532), .B(n260), .CI(n509), .CO(n539), .S(n538) );
  ad01d0 U795 ( .A(n275), .B(n536), .CI(n513), .CO(n543), .S(n542) );
  ad01d0 U796 ( .A(n691), .B(n702), .CI(n693), .CO(n707), .S(n706) );
  ad01d0 U797 ( .A(n482), .B(n484), .CI(n273), .CO(n491), .S(n490) );
  ad01d0 U798 ( .A(n133), .B(n148), .CI(n163), .CO(n379), .S(n378) );
  ad01d0 U799 ( .A(n435), .B(n242), .CI(n107), .CO(n461), .S(n460) );
  ad01d0 U800 ( .A(n121), .B(n151), .CI(n181), .CO(n435), .S(n434) );
  ad01d0 U801 ( .A(n89), .B(n119), .CI(n392), .CO(n399), .S(n398) );
  ad01d0 U802 ( .A(n92), .B(n441), .CI(n460), .CO(n467), .S(n466) );
  ad01d0 U803 ( .A(n91), .B(n419), .CI(n436), .CO(n443), .S(n442) );
  ad01d0 U804 ( .A(n439), .B(n257), .CI(n458), .CO(n465), .S(n464) );
  ad01d0 U805 ( .A(n445), .B(n77), .CI(n464), .CO(n471), .S(n470) );
  ad01d0 U806 ( .A(n469), .B(n78), .CI(n490), .CO(n497), .S(n496) );
  ad01d0 U807 ( .A(n110), .B(n517), .CI(n542), .CO(n549), .S(n548) );
  ad01d0 U808 ( .A(n461), .B(n108), .CI(n463), .CO(n489), .S(n488) );
  ad01d0 U809 ( .A(n376), .B(n365), .CI(n367), .CO(n385), .S(n384) );
  ad01d0 U810 ( .A(n323), .B(n113), .CI(n68), .CO(n329), .S(n328) );
  ad01d0 U811 ( .A(n342), .B(n344), .CI(n339), .CO(n349), .S(n348) );
  ad01d0 U812 ( .A(n347), .B(n356), .CI(n349), .CO(n361), .S(n360) );
  ad01d0 U813 ( .A(n714), .B(n707), .CI(n716), .CO(n719), .S(n718) );
  ad01d0 U814 ( .A(n722), .B(n717), .CI(n724), .CO(n727), .S(n726) );
  ad01d0 U815 ( .A(n75), .B(n414), .CI(n401), .CO(n423), .S(n422) );
  ad01d0 U816 ( .A(n84), .B(n129), .CI(n327), .CO(n335), .S(n334) );
  ad01d0 U817 ( .A(n87), .B(n177), .CI(n362), .CO(n369), .S(n368) );
  ad01d0 U818 ( .A(n122), .B(n227), .CI(n433), .CO(n459), .S(n458) );
  ad01d0 U819 ( .A(n140), .B(n534), .CI(n511), .CO(n541), .S(n540) );
  ad01d0 U820 ( .A(n213), .B(n153), .CI(n183), .CO(n479), .S(n478) );
  ad01d0 U821 ( .A(n216), .B(n201), .CI(n186), .CO(n559), .S(n558) );
  ad01d0 U822 ( .A(n264), .B(n609), .CI(n204), .CO(n633), .S(n632) );
  ad01d0 U823 ( .A(n277), .B(n565), .CI(n157), .CO(n593), .S(n592) );
  ad01d0 U824 ( .A(n278), .B(n589), .CI(n173), .CO(n615), .S(n614) );
  ad01d0 U825 ( .A(n218), .B(n233), .CI(n248), .CO(n609), .S(n608) );
  ad01d0 U826 ( .A(n250), .B(n235), .CI(n265), .CO(n651), .S(n650) );
  ad01d0 U827 ( .A(n190), .B(n652), .CI(n637), .CO(n659), .S(n658) );
  ad01d0 U828 ( .A(n268), .B(n283), .CI(n253), .CO(n699), .S(n698) );
  ad01d0 U829 ( .A(n588), .B(n292), .CI(n567), .CO(n595), .S(n594) );
  ad01d0 U830 ( .A(n559), .B(n247), .CI(n187), .CO(n587), .S(n586) );
  ad01d0 U831 ( .A(n480), .B(n459), .CI(n258), .CO(n487), .S(n486) );
  ad01d0 U832 ( .A(n564), .B(n541), .CI(n291), .CO(n571), .S(n570) );
  ad01d0 U833 ( .A(n610), .B(n591), .CI(n293), .CO(n617), .S(n616) );
  ad01d0 U834 ( .A(n366), .B(n357), .CI(n368), .CO(n373), .S(n372) );
  ad01d0 U835 ( .A(n394), .B(n381), .CI(n383), .CO(n403), .S(n402) );
  ad01d0 U836 ( .A(n471), .B(n492), .CI(n494), .CO(n499), .S(n498) );
  ad01d0 U837 ( .A(n400), .B(n387), .CI(n402), .CO(n407), .S(n406) );
  ad01d0 U838 ( .A(n447), .B(n466), .CI(n468), .CO(n473), .S(n472) );
  ad01d0 U839 ( .A(n425), .B(n442), .CI(n444), .CO(n449), .S(n448) );
  ad01d0 U840 ( .A(n405), .B(n420), .CI(n422), .CO(n427), .S(n426) );
  ad01d0 U841 ( .A(n568), .B(n547), .CI(n570), .CO(n577), .S(n576) );
  ad01d0 U842 ( .A(n574), .B(n553), .CI(n576), .CO(n581), .S(n580) );
  ad01d0 U843 ( .A(n548), .B(n525), .CI(n550), .CO(n555), .S(n554) );
  ad01d0 U844 ( .A(n677), .B(n690), .CI(n679), .CO(n695), .S(n694) );
  ad01d0 U845 ( .A(n661), .B(n676), .CI(n663), .CO(n681), .S(n680) );
  ad01d0 U846 ( .A(n497), .B(n520), .CI(n522), .CO(n527), .S(n526) );
  ad01d0 U847 ( .A(n643), .B(n660), .CI(n645), .CO(n665), .S(n664) );
  ad01d0 U848 ( .A(n703), .B(n712), .CI(n705), .CO(n717), .S(n716) );
  ad01d0 U849 ( .A(n713), .B(n720), .CI(n715), .CO(n725), .S(n724) );
  ad01d0 U850 ( .A(n73), .B(n103), .CI(n178), .CO(n383), .S(n382) );
  ad01d0 U851 ( .A(n125), .B(n538), .CI(n290), .CO(n545), .S(n544) );
  ad01d0 U852 ( .A(n377), .B(n209), .CI(n179), .CO(n397), .S(n396) );
  ad01d0 U853 ( .A(n166), .B(n411), .CI(n211), .CO(n433), .S(n432) );
  ad01d0 U854 ( .A(n72), .B(n147), .CI(n102), .CO(n367), .S(n366) );
  ad01d0 U855 ( .A(n134), .B(n149), .CI(n164), .CO(n395), .S(n394) );
  ad01d0 U856 ( .A(n259), .B(n506), .CI(n124), .CO(n513), .S(n512) );
  ad01d0 U857 ( .A(n537), .B(n560), .CI(n276), .CO(n567), .S(n566) );
  ad01d0 U858 ( .A(n453), .B(n476), .CI(n138), .CO(n481), .S(n480) );
  ad01d0 U859 ( .A(n562), .B(n539), .CI(n141), .CO(n569), .S(n568) );
  ad01d0 U860 ( .A(n199), .B(n477), .CI(n184), .CO(n505), .S(n504) );
  ad01d0 U861 ( .A(n231), .B(n531), .CI(n246), .CO(n561), .S(n560) );
  ad01d0 U862 ( .A(n203), .B(n585), .CI(n263), .CO(n611), .S(n610) );
  ad01d0 U863 ( .A(n137), .B(n167), .CI(n452), .CO(n457), .S(n456) );
  ad01d0 U864 ( .A(n633), .B(n205), .CI(n650), .CO(n655), .S(n654) );
  ad01d0 U865 ( .A(n189), .B(n613), .CI(n632), .CO(n637), .S(n636) );
  ad01d0 U866 ( .A(n672), .B(n659), .CI(n674), .CO(n679), .S(n678) );
  ad01d0 U867 ( .A(n641), .B(n656), .CI(n658), .CO(n663), .S(n662) );
  ad01d0 U868 ( .A(n618), .B(n599), .CI(n620), .CO(n625), .S(n624) );
  ad01d0 U869 ( .A(n575), .B(n596), .CI(n598), .CO(n603), .S(n602) );
  ad01d0 U870 ( .A(n638), .B(n621), .CI(n640), .CO(n645), .S(n644) );
  ad01d0 U871 ( .A(n687), .B(n689), .CI(n700), .CO(n705), .S(n704) );
  ad01d0 U872 ( .A(n686), .B(n675), .CI(n688), .CO(n693), .S(n692) );
  ad01d0 U873 ( .A(n332), .B(n69), .CI(n329), .CO(n337), .S(n336) );
  ad01d0 U874 ( .A(n135), .B(n410), .CI(n395), .CO(n417), .S(n416) );
  ad01d0 U875 ( .A(n228), .B(n455), .CI(n457), .CO(n483), .S(n482) );
  ad01d0 U876 ( .A(n139), .B(n504), .CI(n483), .CO(n511), .S(n510) );
  ad01d0 U877 ( .A(n549), .B(n572), .CI(n551), .CO(n579), .S(n578) );
  ad01d0 U878 ( .A(n738), .B(n737), .CI(n891), .CO(n892), .S(product[29]) );
  ad01d0 U879 ( .A(n723), .B(n725), .CI(n730), .CO(n733), .S(n732) );
  ad01d0 U880 ( .A(n729), .B(n734), .CI(n731), .CO(n737), .S(n736) );
  inv0d1 U881 ( .I(b[13]), .ZN(n61) );
  ad01d0 U882 ( .A(n238), .B(n223), .CI(n698), .CO(n703), .S(n702) );
  ad01d0 U883 ( .A(n684), .B(n207), .CI(n673), .CO(n691), .S(n690) );
  ad01d0 U884 ( .A(n175), .B(n654), .CI(n639), .CO(n661), .S(n660) );
  ad01d0 U885 ( .A(n295), .B(n635), .CI(n310), .CO(n657), .S(n656) );
  ad01d0 U886 ( .A(n191), .B(n670), .CI(n657), .CO(n677), .S(n676) );
  ad01d0 U887 ( .A(n314), .B(n699), .CI(n254), .CO(n713), .S(n712) );
  ad01d0 U888 ( .A(n399), .B(n412), .CI(n240), .CO(n421), .S(n420) );
  ad01d0 U889 ( .A(n192), .B(n117), .CI(n162), .CO(n365), .S(n364) );
  ad01d0 U890 ( .A(n306), .B(n543), .CI(n126), .CO(n573), .S(n572) );
  ad01d0 U891 ( .A(n294), .B(n309), .CI(n615), .CO(n639), .S(n638) );
  ad01d0 U892 ( .A(n612), .B(n308), .CI(n593), .CO(n619), .S(n618) );
  ad01d0 U893 ( .A(n239), .B(n701), .CI(n710), .CO(n715), .S(n714) );
  ad01d0 U894 ( .A(n128), .B(n326), .CI(n325), .CO(n331), .S(n330) );
  ad01d0 U895 ( .A(n71), .B(n176), .CI(n343), .CO(n357), .S(n356) );
  ad01d0 U896 ( .A(n307), .B(n590), .CI(n569), .CO(n597), .S(n596) );
  ad01d0 U897 ( .A(n443), .B(n462), .CI(n272), .CO(n469), .S(n468) );
  ad01d0 U898 ( .A(n566), .B(n111), .CI(n545), .CO(n575), .S(n574) );
  ad01d0 U899 ( .A(n160), .B(n335), .CI(n337), .CO(n347), .S(n346) );
  ad01d0 U900 ( .A(n256), .B(n421), .CI(n76), .CO(n445), .S(n444) );
  ad01d0 U901 ( .A(n118), .B(n363), .CI(n208), .CO(n381), .S(n380) );
  ad01d0 U902 ( .A(n142), .B(n127), .CI(n592), .CO(n599), .S(n598) );
  ad01d0 U903 ( .A(n312), .B(n671), .CI(n222), .CO(n689), .S(n688) );
  ad01d0 U904 ( .A(n158), .B(n143), .CI(n614), .CO(n621), .S(n620) );
  ad01d0 U905 ( .A(n174), .B(n634), .CI(n159), .CO(n641), .S(n640) );
  ad01d0 U906 ( .A(n311), .B(n206), .CI(n655), .CO(n675), .S(n674) );
  ad01d0 U907 ( .A(n298), .B(n685), .CI(n313), .CO(n701), .S(n700) );
  ad01d0 U908 ( .A(n467), .B(n288), .CI(n488), .CO(n495), .S(n494) );
  ad01d0 U909 ( .A(n515), .B(n305), .CI(n540), .CO(n547), .S(n546) );
  ad01d0 U910 ( .A(n514), .B(n493), .CI(n79), .CO(n523), .S(n522) );
  ad01d0 U911 ( .A(n321), .B(n67), .CI(n112), .CO(n325), .S(n324) );
  ad01d0 U912 ( .A(n379), .B(n74), .CI(n224), .CO(n401), .S(n400) );
  ad01d0 U913 ( .A(n491), .B(n304), .CI(n94), .CO(n521), .S(n520) );
  ad01d0 U914 ( .A(n144), .B(n331), .CI(n334), .CO(n339), .S(n338) );
  ad01d0 U915 ( .A(n95), .B(n519), .CI(n521), .CO(n551), .S(n550) );
  ad01d0 U916 ( .A(n285), .B(n300), .CI(n315), .CO(n721), .S(n720) );
  ad01d0 U917 ( .A(n301), .B(n316), .CI(n286), .CO(n729), .S(n728) );
  ad01d0 U918 ( .A(n270), .B(n255), .CI(n711), .CO(n723), .S(n722) );
  ad01d0 U919 ( .A(n271), .B(n721), .CI(n728), .CO(n731), .S(n730) );
  ad01d0 U920 ( .A(n317), .B(n302), .CI(n287), .CO(n735), .S(n734) );
  ad01d0 U921 ( .A(n318), .B(n303), .CI(n735), .CO(n739), .S(n738) );
  inv0d1 U922 ( .I(n767), .ZN(n769) );
  inv0d1 U923 ( .I(b[1]), .ZN(n49) );
  inv0d1 U924 ( .I(a[1]), .ZN(n33) );
  inv0d1 U925 ( .I(a[2]), .ZN(n34) );
  inv0d1 U926 ( .I(b[4]), .ZN(n52) );
  inv0d1 U927 ( .I(a[3]), .ZN(n35) );
  inv0d1 U928 ( .I(a[4]), .ZN(n36) );
  inv0d1 U929 ( .I(b[3]), .ZN(n51) );
  aoi21d1 U930 ( .B1(n960), .B2(n769), .A(n772), .ZN(n774) );
  inv0d1 U931 ( .I(n770), .ZN(n772) );
  aoi21d1 U932 ( .B1(n962), .B2(n777), .A(n780), .ZN(n782) );
  inv0d1 U933 ( .I(n778), .ZN(n780) );
  inv0d1 U934 ( .I(b[2]), .ZN(n50) );
  aoi21d1 U935 ( .B1(n813), .B2(n958), .A(n816), .ZN(n818) );
  inv0d1 U936 ( .I(n814), .ZN(n816) );
  inv0d1 U937 ( .I(n786), .ZN(n788) );
  inv0d1 U938 ( .I(n794), .ZN(n796) );
  inv0d1 U939 ( .I(a[10]), .ZN(n42) );
  inv0d1 U940 ( .I(a[7]), .ZN(n39) );
  inv0d1 U941 ( .I(a[5]), .ZN(n37) );
  inv0d1 U942 ( .I(b[5]), .ZN(n53) );
  inv0d1 U943 ( .I(a[8]), .ZN(n40) );
  inv0d1 U944 ( .I(b[6]), .ZN(n54) );
  inv0d1 U945 ( .I(b[8]), .ZN(n56) );
  inv0d1 U946 ( .I(a[6]), .ZN(n38) );
  inv0d1 U947 ( .I(n886), .ZN(n765) );
  inv0d1 U948 ( .I(a[14]), .ZN(n46) );
  inv0d1 U949 ( .I(a[13]), .ZN(n45) );
  inv0d1 U950 ( .I(a[15]), .ZN(n47) );
  inv0d1 U951 ( .I(b[9]), .ZN(n57) );
  inv0d1 U952 ( .I(a[9]), .ZN(n41) );
  inv0d1 U953 ( .I(n800), .ZN(n748) );
  inv0d1 U954 ( .I(b[7]), .ZN(n55) );
  inv0d1 U955 ( .I(a[11]), .ZN(n43) );
  inv0d1 U956 ( .I(a[12]), .ZN(n44) );
  inv0d1 U957 ( .I(b[15]), .ZN(n63) );
  aoi21d1 U958 ( .B1(n819), .B2(n956), .A(n822), .ZN(n824) );
  inv0d1 U959 ( .I(n820), .ZN(n822) );
  inv0d1 U960 ( .I(n804), .ZN(n749) );
  inv0d1 U961 ( .I(b[10]), .ZN(n58) );
  inv0d1 U962 ( .I(b[12]), .ZN(n60) );
  inv0d1 U963 ( .I(n873), .ZN(n875) );
  inv0d1 U964 ( .I(n812), .ZN(n751) );
  inv0d1 U965 ( .I(n776), .ZN(n742) );
  inv0d1 U966 ( .I(n792), .ZN(n746) );
  inv0d1 U967 ( .I(n825), .ZN(n827) );
  inv0d1 U968 ( .I(n784), .ZN(n744) );
  aoi21d1 U969 ( .B1(n961), .B2(n785), .A(n788), .ZN(n790) );
  aoi21d1 U970 ( .B1(n793), .B2(n959), .A(n796), .ZN(n798) );
  inv0d1 U971 ( .I(n842), .ZN(n844) );
  inv0d1 U972 ( .I(n807), .ZN(n750) );
  inv0d1 U973 ( .I(b[11]), .ZN(n59) );
  inv0d1 U974 ( .I(n864), .ZN(n761) );
  inv0d1 U975 ( .I(n879), .ZN(n764) );
  inv0d1 U976 ( .I(n834), .ZN(n755) );
  inv0d1 U977 ( .I(b[14]), .ZN(n62) );
  inv0d1 U978 ( .I(n869), .ZN(n871) );
  inv0d1 U979 ( .I(n837), .ZN(n756) );
  inv0d1 U980 ( .I(n867), .ZN(n762) );
  inv0d1 U981 ( .I(n853), .ZN(n759) );
  inv0d1 U982 ( .I(n856), .ZN(n760) );
  inv0d1 U983 ( .I(n874), .ZN(n876) );
  inv0d1 U984 ( .I(n868), .ZN(n870) );
  aoi21d1 U985 ( .B1(n868), .B2(n881), .A(n880), .ZN(n882) );
  inv0d1 U986 ( .I(n843), .ZN(n845) );
  aoi21d1 U987 ( .B1(n957), .B2(n822), .A(n827), .ZN(n829) );
  inv0d1 U988 ( .I(n840), .ZN(n841) );
  aoi21d1 U989 ( .B1(n831), .B2(n839), .A(n838), .ZN(n840) );
  inv0d1 U990 ( .I(n848), .ZN(n758) );
  aoi21d1 U991 ( .B1(n841), .B2(n850), .A(n849), .ZN(n851) );
  aoi21d1 U992 ( .B1(n849), .B2(n858), .A(n857), .ZN(n859) );
  inv0d1 U993 ( .I(n861), .ZN(n862) );
  inv0d1 U994 ( .I(a[0]), .ZN(n32) );
  inv0d1 U995 ( .I(b[0]), .ZN(n48) );
  inv0d1 U996 ( .I(n801), .ZN(n802) );
  inv0d1 U997 ( .I(n818), .ZN(n819) );
  inv0d1 U998 ( .I(n831), .ZN(n832) );
  ad01d0 U999 ( .A(n319), .B(n739), .CI(n892), .CO(product[31]), .S(
        product[30]) );
endmodule


module BLENDER_DW_mult_uns_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n742, n744, n746, n748, n749, n750, n751, n755, n756, n758, n759,
         n760, n761, n762, n764, n765, n767, n769, n770, n772, n774, n775,
         n776, n777, n778, n780, n782, n783, n784, n785, n786, n788, n790,
         n791, n792, n793, n794, n796, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n816, n818, n819, n820, n822, n824, n825, n827, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n890, n891, n892, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n956, n957, n958, n959, n960,
         n961, n962, n963, n965, n966, n967;

  nr02d0 U33 ( .A1(n32), .A2(n48), .ZN(product[0]) );
  nr02d0 U34 ( .A1(n49), .A2(n32), .ZN(n65) );
  nr02d0 U35 ( .A1(n50), .A2(n32), .ZN(n66) );
  nr02d0 U36 ( .A1(n51), .A2(n32), .ZN(n67) );
  nr02d0 U37 ( .A1(n52), .A2(n32), .ZN(n68) );
  nr02d0 U38 ( .A1(n53), .A2(n32), .ZN(n69) );
  nr02d0 U39 ( .A1(n54), .A2(n32), .ZN(n70) );
  nr02d0 U40 ( .A1(n55), .A2(n32), .ZN(n71) );
  nr02d0 U41 ( .A1(n56), .A2(n32), .ZN(n72) );
  nr02d0 U42 ( .A1(n57), .A2(n32), .ZN(n73) );
  nr02d0 U43 ( .A1(n58), .A2(n32), .ZN(n74) );
  nr02d0 U44 ( .A1(n59), .A2(n32), .ZN(n75) );
  nr02d0 U45 ( .A1(n60), .A2(n32), .ZN(n76) );
  nr02d0 U46 ( .A1(n61), .A2(n32), .ZN(n77) );
  nr02d0 U47 ( .A1(n62), .A2(n32), .ZN(n78) );
  nr02d0 U48 ( .A1(n63), .A2(n32), .ZN(n79) );
  nr02d0 U49 ( .A1(n33), .A2(n48), .ZN(n80) );
  nr02d0 U50 ( .A1(n49), .A2(n33), .ZN(n81) );
  nr02d0 U51 ( .A1(n50), .A2(n33), .ZN(n82) );
  nr02d0 U52 ( .A1(n51), .A2(n33), .ZN(n83) );
  nr02d0 U53 ( .A1(n52), .A2(n33), .ZN(n84) );
  nr02d0 U54 ( .A1(n53), .A2(n33), .ZN(n85) );
  nr02d0 U55 ( .A1(n54), .A2(n33), .ZN(n86) );
  nr02d0 U56 ( .A1(n55), .A2(n33), .ZN(n87) );
  nr02d0 U57 ( .A1(n56), .A2(n33), .ZN(n88) );
  nr02d0 U58 ( .A1(n57), .A2(n33), .ZN(n89) );
  nr02d0 U59 ( .A1(n58), .A2(n33), .ZN(n90) );
  nr02d0 U60 ( .A1(n59), .A2(n33), .ZN(n91) );
  nr02d0 U61 ( .A1(n60), .A2(n33), .ZN(n92) );
  nr02d0 U62 ( .A1(n61), .A2(n33), .ZN(n93) );
  nr02d0 U63 ( .A1(n62), .A2(n33), .ZN(n94) );
  nr02d0 U64 ( .A1(n63), .A2(n33), .ZN(n95) );
  nr02d0 U65 ( .A1(n34), .A2(n48), .ZN(n96) );
  nr02d0 U66 ( .A1(n34), .A2(n49), .ZN(n97) );
  nr02d0 U67 ( .A1(n50), .A2(n34), .ZN(n98) );
  nr02d0 U68 ( .A1(n51), .A2(n34), .ZN(n99) );
  nr02d0 U69 ( .A1(n52), .A2(n34), .ZN(n100) );
  nr02d0 U70 ( .A1(n53), .A2(n34), .ZN(n101) );
  nr02d0 U71 ( .A1(n54), .A2(n34), .ZN(n102) );
  nr02d0 U72 ( .A1(n55), .A2(n34), .ZN(n103) );
  nr02d0 U73 ( .A1(n56), .A2(n34), .ZN(n104) );
  nr02d0 U74 ( .A1(n57), .A2(n34), .ZN(n105) );
  nr02d0 U75 ( .A1(n58), .A2(n34), .ZN(n106) );
  nr02d0 U76 ( .A1(n59), .A2(n34), .ZN(n107) );
  nr02d0 U77 ( .A1(n60), .A2(n34), .ZN(n108) );
  nr02d0 U78 ( .A1(n61), .A2(n34), .ZN(n109) );
  nr02d0 U79 ( .A1(n62), .A2(n34), .ZN(n110) );
  nr02d0 U80 ( .A1(n63), .A2(n34), .ZN(n111) );
  nr02d0 U81 ( .A1(n35), .A2(n48), .ZN(n112) );
  nr02d0 U82 ( .A1(n35), .A2(n49), .ZN(n113) );
  nr02d0 U83 ( .A1(n35), .A2(n50), .ZN(n114) );
  nr02d0 U84 ( .A1(n51), .A2(n35), .ZN(n115) );
  nr02d0 U85 ( .A1(n52), .A2(n35), .ZN(n116) );
  nr02d0 U86 ( .A1(n53), .A2(n35), .ZN(n117) );
  nr02d0 U87 ( .A1(n54), .A2(n35), .ZN(n118) );
  nr02d0 U88 ( .A1(n55), .A2(n35), .ZN(n119) );
  nr02d0 U89 ( .A1(n56), .A2(n35), .ZN(n120) );
  nr02d0 U90 ( .A1(n57), .A2(n35), .ZN(n121) );
  nr02d0 U91 ( .A1(n58), .A2(n35), .ZN(n122) );
  nr02d0 U92 ( .A1(n59), .A2(n35), .ZN(n123) );
  nr02d0 U93 ( .A1(n60), .A2(n35), .ZN(n124) );
  nr02d0 U94 ( .A1(n61), .A2(n35), .ZN(n125) );
  nr02d0 U95 ( .A1(n62), .A2(n35), .ZN(n126) );
  nr02d0 U96 ( .A1(n63), .A2(n35), .ZN(n127) );
  nr02d0 U97 ( .A1(n36), .A2(n48), .ZN(n128) );
  nr02d0 U98 ( .A1(n36), .A2(n49), .ZN(n129) );
  nr02d0 U99 ( .A1(n36), .A2(n50), .ZN(n130) );
  nr02d0 U100 ( .A1(n51), .A2(n36), .ZN(n131) );
  nr02d0 U101 ( .A1(n52), .A2(n36), .ZN(n132) );
  nr02d0 U102 ( .A1(n53), .A2(n36), .ZN(n133) );
  nr02d0 U103 ( .A1(n54), .A2(n36), .ZN(n134) );
  nr02d0 U104 ( .A1(n55), .A2(n36), .ZN(n135) );
  nr02d0 U105 ( .A1(n56), .A2(n36), .ZN(n136) );
  nr02d0 U106 ( .A1(n57), .A2(n36), .ZN(n137) );
  nr02d0 U107 ( .A1(n58), .A2(n36), .ZN(n138) );
  nr02d0 U108 ( .A1(n59), .A2(n36), .ZN(n139) );
  nr02d0 U109 ( .A1(n60), .A2(n36), .ZN(n140) );
  nr02d0 U110 ( .A1(n61), .A2(n36), .ZN(n141) );
  nr02d0 U111 ( .A1(n62), .A2(n36), .ZN(n142) );
  nr02d0 U112 ( .A1(n63), .A2(n36), .ZN(n143) );
  nr02d0 U113 ( .A1(n37), .A2(n48), .ZN(n144) );
  nr02d0 U114 ( .A1(n37), .A2(n49), .ZN(n145) );
  nr02d0 U115 ( .A1(n37), .A2(n50), .ZN(n146) );
  nr02d0 U116 ( .A1(n37), .A2(n51), .ZN(n147) );
  nr02d0 U117 ( .A1(n37), .A2(n52), .ZN(n148) );
  nr02d0 U118 ( .A1(n53), .A2(n37), .ZN(n149) );
  nr02d0 U119 ( .A1(n54), .A2(n37), .ZN(n150) );
  nr02d0 U120 ( .A1(n55), .A2(n37), .ZN(n151) );
  nr02d0 U121 ( .A1(n56), .A2(n37), .ZN(n152) );
  nr02d0 U122 ( .A1(n57), .A2(n37), .ZN(n153) );
  nr02d0 U123 ( .A1(n58), .A2(n37), .ZN(n154) );
  nr02d0 U124 ( .A1(n59), .A2(n37), .ZN(n155) );
  nr02d0 U125 ( .A1(n60), .A2(n37), .ZN(n156) );
  nr02d0 U126 ( .A1(n61), .A2(n37), .ZN(n157) );
  nr02d0 U127 ( .A1(n62), .A2(n37), .ZN(n158) );
  nr02d0 U128 ( .A1(n63), .A2(n37), .ZN(n159) );
  nr02d0 U129 ( .A1(n38), .A2(n48), .ZN(n160) );
  nr02d0 U130 ( .A1(n38), .A2(n49), .ZN(n161) );
  nr02d0 U131 ( .A1(n38), .A2(n50), .ZN(n162) );
  nr02d0 U132 ( .A1(n38), .A2(n51), .ZN(n163) );
  nr02d0 U133 ( .A1(n38), .A2(n52), .ZN(n164) );
  nr02d0 U134 ( .A1(n53), .A2(n38), .ZN(n165) );
  nr02d0 U135 ( .A1(n54), .A2(n38), .ZN(n166) );
  nr02d0 U136 ( .A1(n55), .A2(n38), .ZN(n167) );
  nr02d0 U137 ( .A1(n56), .A2(n38), .ZN(n168) );
  nr02d0 U138 ( .A1(n57), .A2(n38), .ZN(n169) );
  nr02d0 U139 ( .A1(n58), .A2(n38), .ZN(n170) );
  nr02d0 U140 ( .A1(n59), .A2(n38), .ZN(n171) );
  nr02d0 U141 ( .A1(n60), .A2(n38), .ZN(n172) );
  nr02d0 U142 ( .A1(n61), .A2(n38), .ZN(n173) );
  nr02d0 U143 ( .A1(n62), .A2(n38), .ZN(n174) );
  nr02d0 U144 ( .A1(n63), .A2(n38), .ZN(n175) );
  nr02d0 U145 ( .A1(n39), .A2(n48), .ZN(n176) );
  nr02d0 U146 ( .A1(n39), .A2(n49), .ZN(n177) );
  nr02d0 U147 ( .A1(n39), .A2(n50), .ZN(n178) );
  nr02d0 U148 ( .A1(n39), .A2(n51), .ZN(n179) );
  nr02d0 U149 ( .A1(n39), .A2(n52), .ZN(n180) );
  nr02d0 U150 ( .A1(n39), .A2(n53), .ZN(n181) );
  nr02d0 U151 ( .A1(n39), .A2(n54), .ZN(n182) );
  nr02d0 U152 ( .A1(n55), .A2(n39), .ZN(n183) );
  nr02d0 U153 ( .A1(n39), .A2(n56), .ZN(n184) );
  nr02d0 U154 ( .A1(n57), .A2(n39), .ZN(n185) );
  nr02d0 U155 ( .A1(n58), .A2(n39), .ZN(n186) );
  nr02d0 U156 ( .A1(n59), .A2(n39), .ZN(n187) );
  nr02d0 U157 ( .A1(n60), .A2(n39), .ZN(n188) );
  nr02d0 U158 ( .A1(n61), .A2(n39), .ZN(n189) );
  nr02d0 U159 ( .A1(n62), .A2(n39), .ZN(n190) );
  nr02d0 U160 ( .A1(n63), .A2(n39), .ZN(n191) );
  nr02d0 U161 ( .A1(n40), .A2(n48), .ZN(n192) );
  nr02d0 U162 ( .A1(n40), .A2(n49), .ZN(n193) );
  nr02d0 U163 ( .A1(n40), .A2(n50), .ZN(n194) );
  nr02d0 U164 ( .A1(n40), .A2(n51), .ZN(n195) );
  nr02d0 U165 ( .A1(n40), .A2(n52), .ZN(n196) );
  nr02d0 U166 ( .A1(n53), .A2(n40), .ZN(n197) );
  nr02d0 U167 ( .A1(n54), .A2(n40), .ZN(n198) );
  nr02d0 U168 ( .A1(n55), .A2(n40), .ZN(n199) );
  nr02d0 U169 ( .A1(n56), .A2(n40), .ZN(n200) );
  nr02d0 U170 ( .A1(n57), .A2(n40), .ZN(n201) );
  nr02d0 U171 ( .A1(n58), .A2(n40), .ZN(n202) );
  nr02d0 U172 ( .A1(n59), .A2(n40), .ZN(n203) );
  nr02d0 U173 ( .A1(n60), .A2(n40), .ZN(n204) );
  nr02d0 U174 ( .A1(n61), .A2(n40), .ZN(n205) );
  nr02d0 U175 ( .A1(n62), .A2(n40), .ZN(n206) );
  nr02d0 U176 ( .A1(n63), .A2(n40), .ZN(n207) );
  nr02d0 U177 ( .A1(n41), .A2(n48), .ZN(n208) );
  nr02d0 U178 ( .A1(n41), .A2(n49), .ZN(n209) );
  nr02d0 U179 ( .A1(n41), .A2(n50), .ZN(n210) );
  nr02d0 U180 ( .A1(n41), .A2(n51), .ZN(n211) );
  nr02d0 U181 ( .A1(n41), .A2(n52), .ZN(n212) );
  nr02d0 U182 ( .A1(n41), .A2(n53), .ZN(n213) );
  nr02d0 U183 ( .A1(n41), .A2(n54), .ZN(n214) );
  nr02d0 U184 ( .A1(n55), .A2(n41), .ZN(n215) );
  nr02d0 U185 ( .A1(n41), .A2(n56), .ZN(n216) );
  nr02d0 U186 ( .A1(n57), .A2(n41), .ZN(n217) );
  nr02d0 U187 ( .A1(n58), .A2(n41), .ZN(n218) );
  nr02d0 U188 ( .A1(n59), .A2(n41), .ZN(n219) );
  nr02d0 U189 ( .A1(n60), .A2(n41), .ZN(n220) );
  nr02d0 U190 ( .A1(n61), .A2(n41), .ZN(n221) );
  nr02d0 U191 ( .A1(n62), .A2(n41), .ZN(n222) );
  nr02d0 U192 ( .A1(n63), .A2(n41), .ZN(n223) );
  nr02d0 U193 ( .A1(n42), .A2(n48), .ZN(n224) );
  nr02d0 U194 ( .A1(n42), .A2(n49), .ZN(n225) );
  nr02d0 U195 ( .A1(n42), .A2(n50), .ZN(n226) );
  nr02d0 U196 ( .A1(n42), .A2(n51), .ZN(n227) );
  nr02d0 U197 ( .A1(n42), .A2(n52), .ZN(n228) );
  nr02d0 U198 ( .A1(n42), .A2(n53), .ZN(n229) );
  nr02d0 U199 ( .A1(n42), .A2(n54), .ZN(n230) );
  nr02d0 U200 ( .A1(n42), .A2(n55), .ZN(n231) );
  nr02d0 U201 ( .A1(n42), .A2(n56), .ZN(n232) );
  nr02d0 U202 ( .A1(n42), .A2(n57), .ZN(n233) );
  nr02d0 U203 ( .A1(n58), .A2(n42), .ZN(n234) );
  nr02d0 U204 ( .A1(n59), .A2(n42), .ZN(n235) );
  nr02d0 U205 ( .A1(n60), .A2(n42), .ZN(n236) );
  nr02d0 U206 ( .A1(n61), .A2(n42), .ZN(n237) );
  nr02d0 U207 ( .A1(n62), .A2(n42), .ZN(n238) );
  nr02d0 U208 ( .A1(n63), .A2(n42), .ZN(n239) );
  nr02d0 U209 ( .A1(n43), .A2(n48), .ZN(n240) );
  nr02d0 U210 ( .A1(n43), .A2(n49), .ZN(n241) );
  nr02d0 U211 ( .A1(n43), .A2(n50), .ZN(n242) );
  nr02d0 U212 ( .A1(n43), .A2(n51), .ZN(n243) );
  nr02d0 U213 ( .A1(n43), .A2(n52), .ZN(n244) );
  nr02d0 U214 ( .A1(n43), .A2(n53), .ZN(n245) );
  nr02d0 U215 ( .A1(n43), .A2(n54), .ZN(n246) );
  nr02d0 U216 ( .A1(n43), .A2(n55), .ZN(n247) );
  nr02d0 U217 ( .A1(n43), .A2(n56), .ZN(n248) );
  nr02d0 U218 ( .A1(n43), .A2(n57), .ZN(n249) );
  nr02d0 U219 ( .A1(n43), .A2(n58), .ZN(n250) );
  nr02d0 U220 ( .A1(n59), .A2(n43), .ZN(n251) );
  nr02d0 U221 ( .A1(n60), .A2(n43), .ZN(n252) );
  nr02d0 U222 ( .A1(n61), .A2(n43), .ZN(n253) );
  nr02d0 U223 ( .A1(n62), .A2(n43), .ZN(n254) );
  nr02d0 U224 ( .A1(n63), .A2(n43), .ZN(n255) );
  nr02d0 U225 ( .A1(n44), .A2(n48), .ZN(n256) );
  nr02d0 U226 ( .A1(n44), .A2(n49), .ZN(n257) );
  nr02d0 U227 ( .A1(n44), .A2(n50), .ZN(n258) );
  nr02d0 U228 ( .A1(n44), .A2(n51), .ZN(n259) );
  nr02d0 U229 ( .A1(n44), .A2(n52), .ZN(n260) );
  nr02d0 U230 ( .A1(n44), .A2(n53), .ZN(n261) );
  nr02d0 U231 ( .A1(n44), .A2(n54), .ZN(n262) );
  nr02d0 U232 ( .A1(n44), .A2(n55), .ZN(n263) );
  nr02d0 U233 ( .A1(n44), .A2(n56), .ZN(n264) );
  nr02d0 U234 ( .A1(n44), .A2(n57), .ZN(n265) );
  nr02d0 U235 ( .A1(n44), .A2(n58), .ZN(n266) );
  nr02d0 U236 ( .A1(n44), .A2(n59), .ZN(n267) );
  nr02d0 U237 ( .A1(n60), .A2(n44), .ZN(n268) );
  nr02d0 U238 ( .A1(n61), .A2(n44), .ZN(n269) );
  nr02d0 U239 ( .A1(n62), .A2(n44), .ZN(n270) );
  nr02d0 U240 ( .A1(n63), .A2(n44), .ZN(n271) );
  nr02d0 U241 ( .A1(n45), .A2(n48), .ZN(n272) );
  nr02d0 U242 ( .A1(n45), .A2(n49), .ZN(n273) );
  nr02d0 U243 ( .A1(n45), .A2(n50), .ZN(n274) );
  nr02d0 U244 ( .A1(n45), .A2(n51), .ZN(n275) );
  nr02d0 U245 ( .A1(n45), .A2(n52), .ZN(n276) );
  nr02d0 U246 ( .A1(n45), .A2(n53), .ZN(n277) );
  nr02d0 U247 ( .A1(n45), .A2(n54), .ZN(n278) );
  nr02d0 U248 ( .A1(n45), .A2(n55), .ZN(n279) );
  nr02d0 U249 ( .A1(n45), .A2(n56), .ZN(n280) );
  nr02d0 U250 ( .A1(n45), .A2(n57), .ZN(n281) );
  nr02d0 U251 ( .A1(n45), .A2(n58), .ZN(n282) );
  nr02d0 U252 ( .A1(n45), .A2(n59), .ZN(n283) );
  nr02d0 U253 ( .A1(n45), .A2(n60), .ZN(n284) );
  nr02d0 U254 ( .A1(n61), .A2(n45), .ZN(n285) );
  nr02d0 U255 ( .A1(n62), .A2(n45), .ZN(n286) );
  nr02d0 U256 ( .A1(n63), .A2(n45), .ZN(n287) );
  nr02d0 U257 ( .A1(n46), .A2(n48), .ZN(n288) );
  nr02d0 U258 ( .A1(n46), .A2(n49), .ZN(n289) );
  nr02d0 U259 ( .A1(n46), .A2(n50), .ZN(n290) );
  nr02d0 U260 ( .A1(n46), .A2(n51), .ZN(n291) );
  nr02d0 U261 ( .A1(n46), .A2(n52), .ZN(n292) );
  nr02d0 U262 ( .A1(n46), .A2(n53), .ZN(n293) );
  nr02d0 U263 ( .A1(n46), .A2(n54), .ZN(n294) );
  nr02d0 U264 ( .A1(n46), .A2(n55), .ZN(n295) );
  nr02d0 U265 ( .A1(n46), .A2(n56), .ZN(n296) );
  nr02d0 U266 ( .A1(n46), .A2(n57), .ZN(n297) );
  nr02d0 U267 ( .A1(n46), .A2(n58), .ZN(n298) );
  nr02d0 U268 ( .A1(n46), .A2(n59), .ZN(n299) );
  nr02d0 U269 ( .A1(n46), .A2(n60), .ZN(n300) );
  nr02d0 U270 ( .A1(n46), .A2(n61), .ZN(n301) );
  nr02d0 U271 ( .A1(n62), .A2(n46), .ZN(n302) );
  nr02d0 U272 ( .A1(n63), .A2(n46), .ZN(n303) );
  nr02d0 U273 ( .A1(n47), .A2(n48), .ZN(n304) );
  nr02d0 U274 ( .A1(n47), .A2(n49), .ZN(n305) );
  nr02d0 U275 ( .A1(n47), .A2(n50), .ZN(n306) );
  nr02d0 U276 ( .A1(n47), .A2(n51), .ZN(n307) );
  nr02d0 U277 ( .A1(n47), .A2(n52), .ZN(n308) );
  nr02d0 U278 ( .A1(n47), .A2(n53), .ZN(n309) );
  nr02d0 U279 ( .A1(n47), .A2(n54), .ZN(n310) );
  nr02d0 U280 ( .A1(n47), .A2(n55), .ZN(n311) );
  nr02d0 U281 ( .A1(n47), .A2(n56), .ZN(n312) );
  nr02d0 U282 ( .A1(n47), .A2(n57), .ZN(n313) );
  nr02d0 U283 ( .A1(n47), .A2(n58), .ZN(n314) );
  nr02d0 U284 ( .A1(n47), .A2(n59), .ZN(n315) );
  nr02d0 U285 ( .A1(n47), .A2(n60), .ZN(n316) );
  nr02d0 U286 ( .A1(n47), .A2(n61), .ZN(n317) );
  nr02d0 U287 ( .A1(n62), .A2(n47), .ZN(n318) );
  nr02d0 U288 ( .A1(n63), .A2(n47), .ZN(n319) );
  ah01d0 U289 ( .A(n81), .B(n96), .CO(n321), .S(n320) );
  ah01d0 U290 ( .A(n97), .B(n82), .CO(n323), .S(n322) );
  ah01d0 U292 ( .A(n98), .B(n113), .CO(n327), .S(n326) );
  ah01d0 U295 ( .A(n114), .B(n129), .CO(n333), .S(n332) );
  ah01d0 U299 ( .A(n130), .B(n115), .CO(n341), .S(n340) );
  ah01d0 U304 ( .A(n131), .B(n116), .CO(n351), .S(n350) );
  ah01d0 U310 ( .A(n132), .B(n192), .CO(n363), .S(n362) );
  ah01d0 U317 ( .A(n193), .B(n148), .CO(n377), .S(n376) );
  ah01d0 U325 ( .A(n194), .B(n164), .CO(n393), .S(n392) );
  ah01d0 U334 ( .A(n195), .B(n120), .CO(n411), .S(n410) );
  ah01d0 U344 ( .A(n196), .B(n136), .CO(n431), .S(n430) );
  ah01d0 U355 ( .A(n152), .B(n197), .CO(n453), .S(n452) );
  ah01d0 U367 ( .A(n168), .B(n198), .CO(n477), .S(n476) );
  ah01d0 U380 ( .A(n214), .B(n184), .CO(n503), .S(n502) );
  ah01d0 U394 ( .A(n200), .B(n185), .CO(n531), .S(n530) );
  nd02d1 U499 ( .A1(n65), .A2(n80), .ZN(n767) );
  nd02d1 U505 ( .A1(n320), .A2(n66), .ZN(n770) );
  nd02d1 U508 ( .A1(n960), .A2(n770), .ZN(n895) );
  xn02d1 U512 ( .A1(n895), .A2(n769), .ZN(product[2]) );
  nd02d1 U513 ( .A1(n324), .A2(n322), .ZN(n775) );
  nr02d0 U514 ( .A1(n324), .A2(n322), .ZN(n776) );
  nd02d1 U516 ( .A1(n742), .A2(n775), .ZN(n896) );
  oai21d1 U517 ( .B1(n776), .B2(n774), .A(n775), .ZN(n777) );
  xr02d1 U518 ( .A1(n896), .A2(n774), .Z(product[3]) );
  nd02d1 U519 ( .A1(n330), .A2(n328), .ZN(n778) );
  nd02d1 U522 ( .A1(n962), .A2(n778), .ZN(n897) );
  xn02d1 U526 ( .A1(n897), .A2(n777), .ZN(product[4]) );
  nd02d1 U527 ( .A1(n338), .A2(n336), .ZN(n783) );
  nr02d0 U528 ( .A1(n338), .A2(n336), .ZN(n784) );
  nd02d1 U530 ( .A1(n744), .A2(n783), .ZN(n898) );
  oai21d1 U531 ( .B1(n784), .B2(n782), .A(n783), .ZN(n785) );
  xr02d1 U532 ( .A1(n898), .A2(n782), .Z(product[5]) );
  nd02d1 U533 ( .A1(n348), .A2(n346), .ZN(n786) );
  nd02d1 U536 ( .A1(n961), .A2(n786), .ZN(n899) );
  xn02d1 U540 ( .A1(n899), .A2(n785), .ZN(product[6]) );
  nd02d1 U541 ( .A1(n360), .A2(n358), .ZN(n791) );
  nr02d0 U542 ( .A1(n360), .A2(n358), .ZN(n792) );
  nd02d1 U544 ( .A1(n746), .A2(n791), .ZN(n900) );
  oai21d1 U545 ( .B1(n792), .B2(n790), .A(n791), .ZN(n793) );
  xr02d1 U546 ( .A1(n900), .A2(n790), .Z(product[7]) );
  nd02d1 U547 ( .A1(n374), .A2(n361), .ZN(n794) );
  nd02d1 U550 ( .A1(n959), .A2(n794), .ZN(n901) );
  xn02d1 U554 ( .A1(n901), .A2(n793), .ZN(product[8]) );
  nd02d1 U555 ( .A1(n390), .A2(n375), .ZN(n799) );
  nr02d0 U556 ( .A1(n390), .A2(n375), .ZN(n800) );
  nd02d1 U558 ( .A1(n748), .A2(n799), .ZN(n902) );
  oai21d1 U559 ( .B1(n798), .B2(n800), .A(n799), .ZN(n801) );
  xr02d1 U561 ( .A1(n798), .A2(n902), .Z(product[9]) );
  nd02d1 U562 ( .A1(n408), .A2(n391), .ZN(n803) );
  nr02d0 U563 ( .A1(n408), .A2(n391), .ZN(n804) );
  nd02d1 U565 ( .A1(n749), .A2(n803), .ZN(n903) );
  oai21d1 U566 ( .B1(n802), .B2(n804), .A(n803), .ZN(n805) );
  xr02d1 U567 ( .A1(n802), .A2(n903), .Z(product[10]) );
  nd02d1 U568 ( .A1(n428), .A2(n409), .ZN(n806) );
  nr02d0 U569 ( .A1(n428), .A2(n409), .ZN(n807) );
  nd02d1 U571 ( .A1(n750), .A2(n806), .ZN(n904) );
  oai21d1 U572 ( .B1(n807), .B2(n803), .A(n806), .ZN(n808) );
  nr02d0 U573 ( .A1(n807), .A2(n804), .ZN(n809) );
  xn02d1 U575 ( .A1(n805), .A2(n904), .ZN(product[11]) );
  nd02d1 U576 ( .A1(n450), .A2(n429), .ZN(n811) );
  nr02d0 U577 ( .A1(n450), .A2(n429), .ZN(n812) );
  nd02d1 U579 ( .A1(n751), .A2(n811), .ZN(n905) );
  oai21d1 U580 ( .B1(n810), .B2(n812), .A(n811), .ZN(n813) );
  xr02d1 U581 ( .A1(n810), .A2(n905), .Z(product[12]) );
  nd02d1 U582 ( .A1(n474), .A2(n451), .ZN(n814) );
  nd02d1 U585 ( .A1(n958), .A2(n814), .ZN(n906) );
  xn02d1 U590 ( .A1(n813), .A2(n906), .ZN(product[13]) );
  nd02d1 U591 ( .A1(n500), .A2(n475), .ZN(n820) );
  nd02d1 U594 ( .A1(n956), .A2(n820), .ZN(n907) );
  xn02d1 U598 ( .A1(n819), .A2(n907), .ZN(product[14]) );
  nd02d1 U599 ( .A1(n528), .A2(n501), .ZN(n825) );
  nd02d1 U602 ( .A1(n957), .A2(n825), .ZN(n908) );
  nd02d1 U606 ( .A1(n957), .A2(n956), .ZN(n830) );
  oai21d1 U607 ( .B1(n830), .B2(n818), .A(n829), .ZN(n831) );
  xr02d1 U609 ( .A1(n824), .A2(n908), .Z(product[15]) );
  nd02d1 U610 ( .A1(n556), .A2(n529), .ZN(n833) );
  nr02d0 U611 ( .A1(n556), .A2(n529), .ZN(n834) );
  nd02d1 U613 ( .A1(n755), .A2(n833), .ZN(n909) );
  oai21d1 U614 ( .B1(n832), .B2(n834), .A(n833), .ZN(n835) );
  xr02d1 U615 ( .A1(n832), .A2(n909), .Z(product[16]) );
  nd02d1 U616 ( .A1(n582), .A2(n557), .ZN(n836) );
  nr02d0 U617 ( .A1(n582), .A2(n557), .ZN(n837) );
  nd02d1 U619 ( .A1(n756), .A2(n836), .ZN(n910) );
  oai21d1 U620 ( .B1(n837), .B2(n833), .A(n836), .ZN(n838) );
  nr02d0 U621 ( .A1(n837), .A2(n834), .ZN(n839) );
  xn02d1 U624 ( .A1(n835), .A2(n910), .ZN(product[17]) );
  nd02d1 U625 ( .A1(n606), .A2(n583), .ZN(n842) );
  nr02d0 U626 ( .A1(n606), .A2(n583), .ZN(n843) );
  nd02d1 U628 ( .A1(n845), .A2(n842), .ZN(n911) );
  xn02d1 U632 ( .A1(n841), .A2(n911), .ZN(product[18]) );
  nd02d1 U633 ( .A1(n628), .A2(n607), .ZN(n847) );
  nr02d0 U634 ( .A1(n628), .A2(n607), .ZN(n848) );
  nd02d1 U636 ( .A1(n758), .A2(n847), .ZN(n912) );
  oai21d1 U637 ( .B1(n848), .B2(n842), .A(n847), .ZN(n849) );
  nr02d0 U638 ( .A1(n848), .A2(n843), .ZN(n850) );
  nd02d1 U641 ( .A1(n648), .A2(n629), .ZN(n852) );
  nr02d0 U642 ( .A1(n648), .A2(n629), .ZN(n853) );
  nd02d1 U644 ( .A1(n759), .A2(n852), .ZN(n913) );
  oai21d1 U645 ( .B1(n851), .B2(n853), .A(n852), .ZN(n854) );
  xr02d1 U646 ( .A1(n851), .A2(n913), .Z(product[20]) );
  nd02d1 U647 ( .A1(n666), .A2(n649), .ZN(n855) );
  nr02d0 U648 ( .A1(n666), .A2(n649), .ZN(n856) );
  nd02d1 U650 ( .A1(n760), .A2(n855), .ZN(n914) );
  oai21d1 U651 ( .B1(n856), .B2(n852), .A(n855), .ZN(n857) );
  nr02d0 U652 ( .A1(n853), .A2(n856), .ZN(n858) );
  nd02d1 U654 ( .A1(n850), .A2(n858), .ZN(n860) );
  oai21d1 U655 ( .B1(n840), .B2(n860), .A(n859), .ZN(n861) );
  xn02d1 U657 ( .A1(n854), .A2(n914), .ZN(product[21]) );
  nd02d1 U658 ( .A1(n682), .A2(n667), .ZN(n863) );
  nr02d0 U659 ( .A1(n682), .A2(n667), .ZN(n864) );
  nd02d1 U661 ( .A1(n761), .A2(n863), .ZN(n915) );
  oai21d1 U662 ( .B1(n862), .B2(n864), .A(n863), .ZN(n865) );
  xr02d1 U663 ( .A1(n862), .A2(n915), .Z(product[22]) );
  nd02d1 U664 ( .A1(n696), .A2(n683), .ZN(n866) );
  nr02d0 U665 ( .A1(n696), .A2(n683), .ZN(n867) );
  nd02d1 U667 ( .A1(n762), .A2(n866), .ZN(n916) );
  oai21d1 U668 ( .B1(n867), .B2(n863), .A(n866), .ZN(n868) );
  nr02d0 U669 ( .A1(n864), .A2(n867), .ZN(n869) );
  oai21d1 U672 ( .B1(n862), .B2(n871), .A(n870), .ZN(n872) );
  xn02d1 U673 ( .A1(n865), .A2(n916), .ZN(product[23]) );
  nd02d1 U674 ( .A1(n708), .A2(n697), .ZN(n873) );
  nr02d0 U675 ( .A1(n708), .A2(n697), .ZN(n874) );
  nd02d1 U677 ( .A1(n876), .A2(n873), .ZN(n917) );
  xn02d1 U681 ( .A1(n872), .A2(n917), .ZN(product[24]) );
  nd02d1 U682 ( .A1(n718), .A2(n709), .ZN(n878) );
  nr02d0 U683 ( .A1(n718), .A2(n709), .ZN(n879) );
  nd02d1 U685 ( .A1(n764), .A2(n878), .ZN(n918) );
  oai21d1 U686 ( .B1(n873), .B2(n879), .A(n878), .ZN(n880) );
  nr02d0 U687 ( .A1(n874), .A2(n879), .ZN(n881) );
  nd02d1 U689 ( .A1(n869), .A2(n881), .ZN(n883) );
  oai21d1 U690 ( .B1(n862), .B2(n883), .A(n882), .ZN(n884) );
  nd02d1 U692 ( .A1(n726), .A2(n719), .ZN(n885) );
  nr02d0 U693 ( .A1(n726), .A2(n719), .ZN(n886) );
  nd02d1 U695 ( .A1(n765), .A2(n885), .ZN(n919) );
  oai21d1 U696 ( .B1(n882), .B2(n886), .A(n885), .ZN(n887) );
  nr02d0 U697 ( .A1(n883), .A2(n886), .ZN(n888) );
  xn02d1 U699 ( .A1(n884), .A2(n919), .ZN(product[26]) );
  ad01d0 U708 ( .A(n727), .B(n732), .CI(n967), .CO(n890), .S(product[27]) );
  or02d1 U709 ( .A1(n500), .A2(n475), .Z(n956) );
  or02d1 U710 ( .A1(n528), .A2(n501), .Z(n957) );
  or02d1 U711 ( .A1(n474), .A2(n451), .Z(n958) );
  or02d1 U712 ( .A1(n374), .A2(n361), .Z(n959) );
  or02d1 U713 ( .A1(n320), .A2(n66), .Z(n960) );
  or02d1 U714 ( .A1(n348), .A2(n346), .Z(n961) );
  or02d1 U715 ( .A1(n330), .A2(n328), .Z(n962) );
  or02d1 U716 ( .A1(n65), .A2(n80), .Z(n963) );
  an02d1 U717 ( .A1(n963), .A2(n767), .Z(product[1]) );
  aoi21d1 U718 ( .B1(n809), .B2(n801), .A(n808), .ZN(n810) );
  xn02d1 U719 ( .A1(n965), .A2(n912), .ZN(product[19]) );
  aor21d1 U720 ( .B1(n841), .B2(n845), .A(n844), .Z(n965) );
  xn02d1 U721 ( .A1(n966), .A2(n918), .ZN(product[25]) );
  aor21d1 U722 ( .B1(n872), .B2(n876), .A(n875), .Z(n966) );
  ad01d0 U723 ( .A(n353), .B(n355), .CI(n364), .CO(n371), .S(n370) );
  ad01d0 U724 ( .A(n416), .B(n403), .CI(n418), .CO(n425), .S(n424) );
  ad01d0 U725 ( .A(n511), .B(n536), .CI(n513), .CO(n543), .S(n542) );
  ad01d0 U726 ( .A(n434), .B(n419), .CI(n436), .CO(n443), .S(n442) );
  ad01d0 U727 ( .A(n437), .B(n454), .CI(n456), .CO(n463), .S(n462) );
  ad01d0 U728 ( .A(n423), .B(n438), .CI(n440), .CO(n447), .S(n446) );
  ad01d0 U729 ( .A(n385), .B(n396), .CI(n398), .CO(n405), .S(n404) );
  ad01d0 U730 ( .A(n376), .B(n365), .CI(n367), .CO(n385), .S(n384) );
  ad01d0 U731 ( .A(n503), .B(n530), .CI(n505), .CO(n535), .S(n534) );
  ad01d0 U732 ( .A(n359), .B(n370), .CI(n372), .CO(n375), .S(n374) );
  ad01d0 U733 ( .A(n473), .B(n496), .CI(n498), .CO(n501), .S(n500) );
  ad01d0 U734 ( .A(n407), .B(n424), .CI(n426), .CO(n429), .S(n428) );
  ad01d0 U735 ( .A(n449), .B(n470), .CI(n472), .CO(n475), .S(n474) );
  ad01d0 U736 ( .A(n427), .B(n446), .CI(n448), .CO(n451), .S(n450) );
  ad01d0 U737 ( .A(n555), .B(n578), .CI(n580), .CO(n583), .S(n582) );
  ad01d0 U738 ( .A(n692), .B(n681), .CI(n694), .CO(n697), .S(n696) );
  ad01d0 U739 ( .A(n389), .B(n404), .CI(n406), .CO(n409), .S(n408) );
  ad01d0 U740 ( .A(n527), .B(n552), .CI(n554), .CO(n557), .S(n556) );
  ad01d0 U741 ( .A(n602), .B(n581), .CI(n604), .CO(n607), .S(n606) );
  ad01d0 U742 ( .A(n644), .B(n627), .CI(n646), .CO(n649), .S(n648) );
  ad01d0 U743 ( .A(n678), .B(n665), .CI(n680), .CO(n683), .S(n682) );
  ad01d0 U744 ( .A(n704), .B(n695), .CI(n706), .CO(n709), .S(n708) );
  ad01d0 U745 ( .A(n373), .B(n386), .CI(n388), .CO(n391), .S(n390) );
  ad01d0 U746 ( .A(n499), .B(n524), .CI(n526), .CO(n529), .S(n528) );
  ad01d0 U747 ( .A(n624), .B(n605), .CI(n626), .CO(n629), .S(n628) );
  ad01d0 U748 ( .A(n662), .B(n647), .CI(n664), .CO(n667), .S(n666) );
  ad01d0 U749 ( .A(n382), .B(n371), .CI(n384), .CO(n389), .S(n388) );
  ad01d0 U750 ( .A(n577), .B(n600), .CI(n579), .CO(n605), .S(n604) );
  ad01d0 U751 ( .A(n623), .B(n642), .CI(n625), .CO(n647), .S(n646) );
  ad01d0 U752 ( .A(n601), .B(n622), .CI(n603), .CO(n627), .S(n626) );
  ad01d0 U753 ( .A(n542), .B(n519), .CI(n544), .CO(n551), .S(n550) );
  aor21d1 U754 ( .B1(n861), .B2(n888), .A(n887), .Z(n967) );
  ad01d0 U755 ( .A(n736), .B(n733), .CI(n890), .CO(n891), .S(product[28]) );
  ad01d0 U756 ( .A(n393), .B(n180), .CI(n105), .CO(n415), .S(n414) );
  ad01d0 U757 ( .A(n215), .B(n230), .CI(n170), .CO(n533), .S(n532) );
  ad01d0 U758 ( .A(n284), .B(n269), .CI(n299), .CO(n711), .S(n710) );
  ad01d0 U759 ( .A(n341), .B(n146), .CI(n161), .CO(n353), .S(n352) );
  ad01d0 U760 ( .A(n243), .B(n123), .CI(n478), .CO(n485), .S(n484) );
  ad01d0 U761 ( .A(n229), .B(n154), .CI(n502), .CO(n507), .S(n506) );
  ad01d0 U762 ( .A(n532), .B(n260), .CI(n509), .CO(n539), .S(n538) );
  ad01d0 U763 ( .A(n245), .B(n155), .CI(n507), .CO(n537), .S(n536) );
  ad01d0 U764 ( .A(n172), .B(n563), .CI(n586), .CO(n591), .S(n590) );
  ad01d0 U765 ( .A(n183), .B(n476), .CI(n228), .CO(n481), .S(n480) );
  ad01d0 U766 ( .A(n630), .B(n279), .CI(n611), .CO(n635), .S(n634) );
  ad01d0 U767 ( .A(n281), .B(n651), .CI(n221), .CO(n671), .S(n670) );
  ad01d0 U768 ( .A(n495), .B(n516), .CI(n518), .CO(n525), .S(n524) );
  ad01d0 U769 ( .A(n595), .B(n597), .CI(n616), .CO(n623), .S(n622) );
  ad01d0 U770 ( .A(n571), .B(n573), .CI(n594), .CO(n601), .S(n600) );
  ad01d0 U771 ( .A(n617), .B(n636), .CI(n619), .CO(n643), .S(n642) );
  ad01d0 U772 ( .A(n100), .B(n333), .CI(n145), .CO(n343), .S(n342) );
  ad01d0 U773 ( .A(n413), .B(n415), .CI(n241), .CO(n439), .S(n438) );
  ad01d0 U774 ( .A(n489), .B(n512), .CI(n289), .CO(n519), .S(n518) );
  ad01d0 U775 ( .A(n212), .B(n182), .CI(n137), .CO(n455), .S(n454) );
  ad01d0 U776 ( .A(n147), .B(n351), .CI(n117), .CO(n365), .S(n364) );
  ad01d0 U777 ( .A(n535), .B(n261), .CI(n156), .CO(n565), .S(n564) );
  ad01d0 U778 ( .A(n268), .B(n283), .CI(n253), .CO(n699), .S(n698) );
  ad01d0 U779 ( .A(n217), .B(n232), .CI(n202), .CO(n585), .S(n584) );
  ad01d0 U780 ( .A(n186), .B(n531), .CI(n246), .CO(n561), .S(n560) );
  ad01d0 U781 ( .A(n234), .B(n249), .CI(n219), .CO(n631), .S(n630) );
  ad01d0 U782 ( .A(n584), .B(n262), .CI(n561), .CO(n589), .S(n588) );
  ad01d0 U783 ( .A(n251), .B(n266), .CI(n236), .CO(n669), .S(n668) );
  ad01d0 U784 ( .A(n631), .B(n220), .CI(n280), .CO(n653), .S(n652) );
  ad01d0 U785 ( .A(n668), .B(n296), .CI(n653), .CO(n673), .S(n672) );
  ad01d0 U786 ( .A(n669), .B(n237), .CI(n297), .CO(n687), .S(n686) );
  ad01d0 U787 ( .A(n179), .B(n119), .CI(n392), .CO(n399), .S(n398) );
  ad01d0 U788 ( .A(n101), .B(n86), .CI(n350), .CO(n355), .S(n354) );
  ad01d0 U789 ( .A(n378), .B(n369), .CI(n380), .CO(n387), .S(n386) );
  ad01d0 U790 ( .A(n465), .B(n93), .CI(n486), .CO(n493), .S(n492) );
  ad01d0 U791 ( .A(n171), .B(n533), .CI(n558), .CO(n563), .S(n562) );
  ad01d0 U792 ( .A(n587), .B(n188), .CI(n608), .CO(n613), .S(n612) );
  ad01d0 U793 ( .A(n487), .B(n109), .CI(n510), .CO(n517), .S(n516) );
  ad01d0 U794 ( .A(n521), .B(n523), .CI(n546), .CO(n553), .S(n552) );
  ad01d0 U795 ( .A(n68), .B(n326), .CI(n325), .CO(n331), .S(n330) );
  ad01d0 U796 ( .A(n395), .B(n90), .CI(n397), .CO(n419), .S(n418) );
  ad01d0 U797 ( .A(n691), .B(n702), .CI(n693), .CO(n707), .S(n706) );
  ad01d0 U798 ( .A(n417), .B(n432), .CI(n91), .CO(n441), .S(n440) );
  ad01d0 U799 ( .A(n135), .B(n410), .CI(n225), .CO(n417), .S(n416) );
  ad01d0 U800 ( .A(n435), .B(n242), .CI(n107), .CO(n461), .S(n460) );
  ad01d0 U801 ( .A(n430), .B(n226), .CI(n106), .CO(n437), .S(n436) );
  ad01d0 U802 ( .A(n463), .B(n484), .CI(n273), .CO(n491), .S(n490) );
  ad01d0 U803 ( .A(n104), .B(n149), .CI(n134), .CO(n395), .S(n394) );
  ad01d0 U804 ( .A(n163), .B(n88), .CI(n118), .CO(n379), .S(n378) );
  ad01d0 U805 ( .A(n165), .B(n150), .CI(n210), .CO(n413), .S(n412) );
  ad01d0 U806 ( .A(n411), .B(n121), .CI(n151), .CO(n435), .S(n434) );
  ad01d0 U807 ( .A(n481), .B(n504), .CI(n259), .CO(n511), .S(n510) );
  ad01d0 U808 ( .A(n213), .B(n153), .CI(n453), .CO(n479), .S(n478) );
  ad01d0 U809 ( .A(n441), .B(n92), .CI(n460), .CO(n467), .S(n466) );
  ad01d0 U810 ( .A(n461), .B(n108), .CI(n482), .CO(n489), .S(n488) );
  ad01d0 U811 ( .A(n345), .B(n352), .CI(n354), .CO(n359), .S(n358) );
  ad01d0 U812 ( .A(n257), .B(n439), .CI(n458), .CO(n465), .S(n464) );
  ad01d0 U813 ( .A(n445), .B(n77), .CI(n464), .CO(n471), .S(n470) );
  ad01d0 U814 ( .A(n469), .B(n78), .CI(n490), .CO(n497), .S(n496) );
  ad01d0 U815 ( .A(n138), .B(n455), .CI(n457), .CO(n483), .S(n482) );
  ad01d0 U816 ( .A(n227), .B(n122), .CI(n433), .CO(n459), .S(n458) );
  ad01d0 U817 ( .A(n85), .B(n335), .CI(n337), .CO(n347), .S(n346) );
  ad01d0 U818 ( .A(n342), .B(n344), .CI(n339), .CO(n349), .S(n348) );
  ad01d0 U819 ( .A(n347), .B(n356), .CI(n349), .CO(n361), .S(n360) );
  ad01d0 U820 ( .A(n714), .B(n707), .CI(n716), .CO(n719), .S(n718) );
  ad01d0 U821 ( .A(n722), .B(n717), .CI(n724), .CO(n727), .S(n726) );
  ad01d0 U822 ( .A(n75), .B(n401), .CI(n414), .CO(n423), .S(n422) );
  ad01d0 U823 ( .A(n99), .B(n84), .CI(n327), .CO(n335), .S(n334) );
  ad01d0 U824 ( .A(n177), .B(n362), .CI(n87), .CO(n369), .S(n368) );
  ad01d0 U825 ( .A(n140), .B(n534), .CI(n275), .CO(n541), .S(n540) );
  ad01d0 U826 ( .A(n125), .B(n538), .CI(n290), .CO(n545), .S(n544) );
  ad01d0 U827 ( .A(n216), .B(n201), .CI(n231), .CO(n559), .S(n558) );
  ad01d0 U828 ( .A(n264), .B(n609), .CI(n204), .CO(n633), .S(n632) );
  ad01d0 U829 ( .A(n278), .B(n589), .CI(n173), .CO(n615), .S(n614) );
  ad01d0 U830 ( .A(n277), .B(n565), .CI(n157), .CO(n593), .S(n592) );
  ad01d0 U831 ( .A(n233), .B(n218), .CI(n248), .CO(n609), .S(n608) );
  ad01d0 U832 ( .A(n247), .B(n559), .CI(n187), .CO(n587), .S(n586) );
  ad01d0 U833 ( .A(n250), .B(n235), .CI(n265), .CO(n651), .S(n650) );
  ad01d0 U834 ( .A(n267), .B(n252), .CI(n282), .CO(n685), .S(n684) );
  ad01d0 U835 ( .A(n564), .B(n291), .CI(n541), .CO(n571), .S(n570) );
  ad01d0 U836 ( .A(n588), .B(n292), .CI(n567), .CO(n595), .S(n594) );
  ad01d0 U837 ( .A(n652), .B(n190), .CI(n637), .CO(n659), .S(n658) );
  ad01d0 U838 ( .A(n459), .B(n480), .CI(n258), .CO(n487), .S(n486) );
  ad01d0 U839 ( .A(n485), .B(n508), .CI(n274), .CO(n515), .S(n514) );
  ad01d0 U840 ( .A(n560), .B(n537), .CI(n276), .CO(n567), .S(n566) );
  ad01d0 U841 ( .A(n610), .B(n591), .CI(n293), .CO(n617), .S(n616) );
  ad01d0 U842 ( .A(n366), .B(n357), .CI(n368), .CO(n373), .S(n372) );
  ad01d0 U843 ( .A(n381), .B(n394), .CI(n383), .CO(n403), .S(n402) );
  ad01d0 U844 ( .A(n471), .B(n492), .CI(n494), .CO(n499), .S(n498) );
  ad01d0 U845 ( .A(n400), .B(n387), .CI(n402), .CO(n407), .S(n406) );
  ad01d0 U846 ( .A(n447), .B(n466), .CI(n468), .CO(n473), .S(n472) );
  ad01d0 U847 ( .A(n425), .B(n442), .CI(n444), .CO(n449), .S(n448) );
  ad01d0 U848 ( .A(n405), .B(n420), .CI(n422), .CO(n427), .S(n426) );
  ad01d0 U849 ( .A(n568), .B(n547), .CI(n570), .CO(n577), .S(n576) );
  ad01d0 U850 ( .A(n574), .B(n553), .CI(n576), .CO(n581), .S(n580) );
  ad01d0 U851 ( .A(n548), .B(n525), .CI(n550), .CO(n555), .S(n554) );
  ad01d0 U852 ( .A(n677), .B(n690), .CI(n679), .CO(n695), .S(n694) );
  ad01d0 U853 ( .A(n661), .B(n676), .CI(n663), .CO(n681), .S(n680) );
  ad01d0 U854 ( .A(n497), .B(n520), .CI(n522), .CO(n527), .S(n526) );
  ad01d0 U855 ( .A(n643), .B(n660), .CI(n645), .CO(n665), .S(n664) );
  ad01d0 U856 ( .A(n703), .B(n712), .CI(n705), .CO(n717), .S(n716) );
  ad01d0 U857 ( .A(n713), .B(n720), .CI(n715), .CO(n725), .S(n724) );
  ad01d0 U858 ( .A(n209), .B(n377), .CI(n89), .CO(n397), .S(n396) );
  ad01d0 U859 ( .A(n178), .B(n73), .CI(n103), .CO(n383), .S(n382) );
  ad01d0 U860 ( .A(n162), .B(n72), .CI(n102), .CO(n367), .S(n366) );
  ad01d0 U861 ( .A(n479), .B(n244), .CI(n139), .CO(n509), .S(n508) );
  ad01d0 U862 ( .A(n483), .B(n506), .CI(n124), .CO(n513), .S(n512) );
  ad01d0 U863 ( .A(n562), .B(n539), .CI(n141), .CO(n569), .S(n568) );
  ad01d0 U864 ( .A(n169), .B(n477), .CI(n199), .CO(n505), .S(n504) );
  ad01d0 U865 ( .A(n166), .B(n211), .CI(n181), .CO(n433), .S(n432) );
  ad01d0 U866 ( .A(n203), .B(n585), .CI(n263), .CO(n611), .S(n610) );
  ad01d0 U867 ( .A(n431), .B(n167), .CI(n452), .CO(n457), .S(n456) );
  ad01d0 U868 ( .A(n329), .B(n331), .CI(n334), .CO(n339), .S(n338) );
  ad01d0 U869 ( .A(n633), .B(n205), .CI(n650), .CO(n655), .S(n654) );
  ad01d0 U870 ( .A(n189), .B(n613), .CI(n632), .CO(n637), .S(n636) );
  ad01d0 U871 ( .A(n672), .B(n659), .CI(n674), .CO(n679), .S(n678) );
  ad01d0 U872 ( .A(n656), .B(n641), .CI(n658), .CO(n663), .S(n662) );
  ad01d0 U873 ( .A(n618), .B(n599), .CI(n620), .CO(n625), .S(n624) );
  ad01d0 U874 ( .A(n596), .B(n575), .CI(n598), .CO(n603), .S(n602) );
  ad01d0 U875 ( .A(n638), .B(n621), .CI(n640), .CO(n645), .S(n644) );
  ad01d0 U876 ( .A(n698), .B(n689), .CI(n700), .CO(n705), .S(n704) );
  ad01d0 U877 ( .A(n686), .B(n675), .CI(n688), .CO(n693), .S(n692) );
  ad01d0 U878 ( .A(n549), .B(n572), .CI(n551), .CO(n579), .S(n578) );
  ad01d0 U879 ( .A(n738), .B(n737), .CI(n891), .CO(n892), .S(product[29]) );
  ad01d0 U880 ( .A(n723), .B(n725), .CI(n730), .CO(n733), .S(n732) );
  ad01d0 U881 ( .A(n729), .B(n734), .CI(n731), .CO(n737), .S(n736) );
  ad01d0 U882 ( .A(n160), .B(n340), .CI(n70), .CO(n345), .S(n344) );
  inv0d1 U883 ( .I(b[12]), .ZN(n60) );
  inv0d1 U884 ( .I(b[13]), .ZN(n61) );
  ad01d0 U885 ( .A(n222), .B(n207), .CI(n673), .CO(n691), .S(n690) );
  ad01d0 U886 ( .A(n238), .B(n223), .CI(n687), .CO(n703), .S(n702) );
  ad01d0 U887 ( .A(n491), .B(n304), .CI(n514), .CO(n521), .S(n520) );
  ad01d0 U888 ( .A(n175), .B(n654), .CI(n639), .CO(n661), .S(n660) );
  ad01d0 U889 ( .A(n191), .B(n670), .CI(n657), .CO(n677), .S(n676) );
  ad01d0 U890 ( .A(n314), .B(n699), .CI(n254), .CO(n713), .S(n712) );
  ad01d0 U891 ( .A(n412), .B(n399), .CI(n240), .CO(n421), .S(n420) );
  ad01d0 U892 ( .A(n176), .B(n343), .CI(n71), .CO(n357), .S(n356) );
  ad01d0 U893 ( .A(n379), .B(n224), .CI(n74), .CO(n401), .S(n400) );
  ad01d0 U894 ( .A(n294), .B(n309), .CI(n615), .CO(n639), .S(n638) );
  ad01d0 U895 ( .A(n612), .B(n308), .CI(n593), .CO(n619), .S(n618) );
  ad01d0 U896 ( .A(n295), .B(n635), .CI(n310), .CO(n657), .S(n656) );
  ad01d0 U897 ( .A(n239), .B(n701), .CI(n710), .CO(n715), .S(n714) );
  ad01d0 U898 ( .A(n306), .B(n543), .CI(n566), .CO(n573), .S(n572) );
  ad01d0 U899 ( .A(n126), .B(n111), .CI(n545), .CO(n575), .S(n574) );
  ad01d0 U900 ( .A(n307), .B(n590), .CI(n569), .CO(n597), .S(n596) );
  ad01d0 U901 ( .A(n110), .B(n517), .CI(n95), .CO(n549), .S(n548) );
  ad01d0 U902 ( .A(n443), .B(n272), .CI(n462), .CO(n469), .S(n468) );
  ad01d0 U903 ( .A(n323), .B(n128), .CI(n83), .CO(n329), .S(n328) );
  ad01d0 U904 ( .A(n256), .B(n421), .CI(n76), .CO(n445), .S(n444) );
  ad01d0 U905 ( .A(n94), .B(n493), .CI(n79), .CO(n523), .S(n522) );
  ad01d0 U906 ( .A(n133), .B(n363), .CI(n208), .CO(n381), .S(n380) );
  ad01d0 U907 ( .A(n142), .B(n127), .CI(n592), .CO(n599), .S(n598) );
  ad01d0 U908 ( .A(n174), .B(n634), .CI(n159), .CO(n641), .S(n640) );
  ad01d0 U909 ( .A(n158), .B(n143), .CI(n614), .CO(n621), .S(n620) );
  ad01d0 U910 ( .A(n312), .B(n671), .CI(n684), .CO(n689), .S(n688) );
  ad01d0 U911 ( .A(n311), .B(n206), .CI(n655), .CO(n675), .S(n674) );
  ad01d0 U912 ( .A(n298), .B(n685), .CI(n313), .CO(n701), .S(n700) );
  ad01d0 U913 ( .A(n467), .B(n288), .CI(n488), .CO(n495), .S(n494) );
  ad01d0 U914 ( .A(n515), .B(n305), .CI(n540), .CO(n547), .S(n546) );
  ad01d0 U915 ( .A(n321), .B(n112), .CI(n67), .CO(n325), .S(n324) );
  ad01d0 U916 ( .A(n144), .B(n332), .CI(n69), .CO(n337), .S(n336) );
  ad01d0 U917 ( .A(n285), .B(n300), .CI(n315), .CO(n721), .S(n720) );
  ad01d0 U918 ( .A(n301), .B(n316), .CI(n286), .CO(n729), .S(n728) );
  ad01d0 U919 ( .A(n270), .B(n255), .CI(n711), .CO(n723), .S(n722) );
  ad01d0 U920 ( .A(n271), .B(n721), .CI(n728), .CO(n731), .S(n730) );
  ad01d0 U921 ( .A(n317), .B(n302), .CI(n287), .CO(n735), .S(n734) );
  ad01d0 U922 ( .A(n318), .B(n303), .CI(n735), .CO(n739), .S(n738) );
  inv0d1 U923 ( .I(a[0]), .ZN(n32) );
  inv0d1 U924 ( .I(n767), .ZN(n769) );
  inv0d1 U925 ( .I(b[1]), .ZN(n49) );
  inv0d1 U926 ( .I(a[1]), .ZN(n33) );
  inv0d1 U927 ( .I(b[2]), .ZN(n50) );
  inv0d1 U928 ( .I(a[4]), .ZN(n36) );
  inv0d1 U929 ( .I(b[4]), .ZN(n52) );
  inv0d1 U930 ( .I(b[3]), .ZN(n51) );
  aoi21d1 U931 ( .B1(n960), .B2(n769), .A(n772), .ZN(n774) );
  inv0d1 U932 ( .I(n770), .ZN(n772) );
  inv0d1 U933 ( .I(a[2]), .ZN(n34) );
  aoi21d1 U934 ( .B1(n813), .B2(n958), .A(n816), .ZN(n818) );
  inv0d1 U935 ( .I(n814), .ZN(n816) );
  inv0d1 U936 ( .I(a[15]), .ZN(n47) );
  inv0d1 U937 ( .I(a[5]), .ZN(n37) );
  inv0d1 U938 ( .I(n778), .ZN(n780) );
  inv0d1 U939 ( .I(b[8]), .ZN(n56) );
  inv0d1 U940 ( .I(a[6]), .ZN(n38) );
  inv0d1 U941 ( .I(b[10]), .ZN(n58) );
  inv0d1 U942 ( .I(n794), .ZN(n796) );
  aoi21d1 U943 ( .B1(n961), .B2(n785), .A(n788), .ZN(n790) );
  inv0d1 U944 ( .I(n786), .ZN(n788) );
  inv0d1 U945 ( .I(a[13]), .ZN(n45) );
  inv0d1 U946 ( .I(b[5]), .ZN(n53) );
  inv0d1 U947 ( .I(n886), .ZN(n765) );
  inv0d1 U948 ( .I(b[7]), .ZN(n55) );
  inv0d1 U949 ( .I(a[9]), .ZN(n41) );
  inv0d1 U950 ( .I(a[14]), .ZN(n46) );
  inv0d1 U951 ( .I(b[6]), .ZN(n54) );
  inv0d1 U952 ( .I(a[10]), .ZN(n42) );
  inv0d1 U953 ( .I(a[11]), .ZN(n43) );
  inv0d1 U954 ( .I(a[12]), .ZN(n44) );
  inv0d1 U955 ( .I(b[9]), .ZN(n57) );
  inv0d1 U956 ( .I(a[7]), .ZN(n39) );
  inv0d1 U957 ( .I(b[14]), .ZN(n62) );
  aoi21d1 U958 ( .B1(n819), .B2(n956), .A(n822), .ZN(n824) );
  inv0d1 U959 ( .I(n820), .ZN(n822) );
  inv0d1 U960 ( .I(n873), .ZN(n875) );
  inv0d1 U961 ( .I(b[15]), .ZN(n63) );
  inv0d1 U962 ( .I(n776), .ZN(n742) );
  inv0d1 U963 ( .I(a[3]), .ZN(n35) );
  inv0d1 U964 ( .I(n792), .ZN(n746) );
  inv0d1 U965 ( .I(n784), .ZN(n744) );
  inv0d1 U966 ( .I(n825), .ZN(n827) );
  inv0d1 U967 ( .I(n800), .ZN(n748) );
  aoi21d1 U968 ( .B1(n962), .B2(n777), .A(n780), .ZN(n782) );
  inv0d1 U969 ( .I(n864), .ZN(n761) );
  inv0d1 U970 ( .I(n812), .ZN(n751) );
  inv0d1 U971 ( .I(n804), .ZN(n749) );
  aoi21d1 U972 ( .B1(n793), .B2(n959), .A(n796), .ZN(n798) );
  inv0d1 U973 ( .I(a[8]), .ZN(n40) );
  inv0d1 U974 ( .I(n842), .ZN(n844) );
  inv0d1 U975 ( .I(n879), .ZN(n764) );
  inv0d1 U976 ( .I(n834), .ZN(n755) );
  inv0d1 U977 ( .I(n807), .ZN(n750) );
  inv0d1 U978 ( .I(b[11]), .ZN(n59) );
  inv0d1 U979 ( .I(n869), .ZN(n871) );
  inv0d1 U980 ( .I(n837), .ZN(n756) );
  inv0d1 U981 ( .I(n867), .ZN(n762) );
  inv0d1 U982 ( .I(n856), .ZN(n760) );
  inv0d1 U983 ( .I(n853), .ZN(n759) );
  inv0d1 U984 ( .I(n874), .ZN(n876) );
  inv0d1 U985 ( .I(n843), .ZN(n845) );
  inv0d1 U986 ( .I(n868), .ZN(n870) );
  aoi21d1 U987 ( .B1(n868), .B2(n881), .A(n880), .ZN(n882) );
  aoi21d1 U988 ( .B1(n957), .B2(n822), .A(n827), .ZN(n829) );
  inv0d1 U989 ( .I(n840), .ZN(n841) );
  aoi21d1 U990 ( .B1(n831), .B2(n839), .A(n838), .ZN(n840) );
  inv0d1 U991 ( .I(n848), .ZN(n758) );
  aoi21d1 U992 ( .B1(n841), .B2(n850), .A(n849), .ZN(n851) );
  aoi21d1 U993 ( .B1(n849), .B2(n858), .A(n857), .ZN(n859) );
  inv0d1 U994 ( .I(n861), .ZN(n862) );
  inv0d1 U995 ( .I(b[0]), .ZN(n48) );
  inv0d1 U996 ( .I(n801), .ZN(n802) );
  inv0d1 U997 ( .I(n818), .ZN(n819) );
  inv0d1 U998 ( .I(n831), .ZN(n832) );
  ad01d0 U999 ( .A(n319), .B(n739), .CI(n892), .CO(product[31]), .S(
        product[30]) );
endmodule


module BLENDER_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n140;

  nr02d0 U17 ( .A1(n17), .A2(A[0]), .ZN(n43) );
  xn02d1 U18 ( .A1(n17), .A2(A[0]), .ZN(DIFF[0]) );
  nd02d1 U19 ( .A1(n18), .A2(A[1]), .ZN(n44) );
  nr02d0 U20 ( .A1(n18), .A2(A[1]), .ZN(n45) );
  nd02d1 U22 ( .A1(n33), .A2(n44), .ZN(n91) );
  oai21d1 U23 ( .B1(n45), .B2(n43), .A(n44), .ZN(n46) );
  xr02d1 U25 ( .A1(n91), .A2(n43), .Z(DIFF[1]) );
  nd02d1 U26 ( .A1(n19), .A2(A[2]), .ZN(n48) );
  nd02d1 U29 ( .A1(n34), .A2(n48), .ZN(n92) );
  oai21d1 U30 ( .B1(n47), .B2(n49), .A(n48), .ZN(n50) );
  xr02d1 U31 ( .A1(n47), .A2(n92), .Z(DIFF[2]) );
  nd02d1 U32 ( .A1(n20), .A2(A[3]), .ZN(n51) );
  nd02d1 U35 ( .A1(n35), .A2(n51), .ZN(n93) );
  oai21d1 U36 ( .B1(n52), .B2(n48), .A(n51), .ZN(n53) );
  nr02d0 U37 ( .A1(n49), .A2(n52), .ZN(n54) );
  xn02d1 U40 ( .A1(n50), .A2(n93), .ZN(DIFF[3]) );
  nd02d1 U41 ( .A1(n21), .A2(A[4]), .ZN(n57) );
  nd02d1 U44 ( .A1(n36), .A2(n57), .ZN(n94) );
  xn02d1 U48 ( .A1(n56), .A2(n94), .ZN(DIFF[4]) );
  nd02d1 U49 ( .A1(n22), .A2(A[5]), .ZN(n62) );
  nd02d1 U52 ( .A1(n37), .A2(n62), .ZN(n95) );
  oai21d1 U53 ( .B1(n63), .B2(n57), .A(n62), .ZN(n64) );
  xr02d1 U56 ( .A1(n61), .A2(n95), .Z(DIFF[5]) );
  nd02d1 U57 ( .A1(n23), .A2(A[6]), .ZN(n67) );
  nd02d1 U60 ( .A1(n38), .A2(n67), .ZN(n96) );
  oai21d1 U61 ( .B1(n66), .B2(n68), .A(n67), .ZN(n69) );
  xr02d1 U62 ( .A1(n66), .A2(n96), .Z(DIFF[6]) );
  nd02d1 U63 ( .A1(n24), .A2(A[7]), .ZN(n70) );
  nd02d1 U66 ( .A1(n39), .A2(n70), .ZN(n97) );
  oai21d1 U67 ( .B1(n71), .B2(n67), .A(n70), .ZN(n72) );
  nr02d0 U68 ( .A1(n68), .A2(n71), .ZN(n73) );
  nd02d1 U70 ( .A1(n65), .A2(n73), .ZN(n75) );
  oai21d1 U71 ( .B1(n55), .B2(n75), .A(n74), .ZN(n76) );
  xn02d1 U73 ( .A1(n69), .A2(n97), .ZN(DIFF[7]) );
  nd02d1 U74 ( .A1(n25), .A2(A[8]), .ZN(n78) );
  nr02d0 U75 ( .A1(n25), .A2(A[8]), .ZN(n79) );
  nd02d1 U77 ( .A1(n40), .A2(n78), .ZN(n98) );
  oai21d1 U78 ( .B1(n77), .B2(n79), .A(n78), .ZN(n80) );
  xr02d1 U79 ( .A1(n77), .A2(n98), .Z(DIFF[8]) );
  nd02d1 U80 ( .A1(n26), .A2(A[9]), .ZN(n81) );
  nr02d0 U81 ( .A1(n26), .A2(A[9]), .ZN(n82) );
  nd02d1 U83 ( .A1(n41), .A2(n81), .ZN(n99) );
  oai21d1 U84 ( .B1(n82), .B2(n78), .A(n81), .ZN(n83) );
  nr02d0 U85 ( .A1(n79), .A2(n82), .ZN(n84) );
  xn02d1 U87 ( .A1(n80), .A2(n99), .ZN(DIFF[9]) );
  xr02d1 U99 ( .A1(n90), .A2(n100), .Z(DIFF[15]) );
  xn02d1 U100 ( .A1(B[15]), .A2(A[15]), .ZN(n100) );
  aor21d1 U101 ( .B1(n76), .B2(n84), .A(n83), .Z(n140) );
  nr02d0 U102 ( .A1(n24), .A2(A[7]), .ZN(n71) );
  nr02d0 U103 ( .A1(n20), .A2(A[3]), .ZN(n52) );
  nr02d0 U104 ( .A1(n22), .A2(A[5]), .ZN(n63) );
  ad01d0 U105 ( .A(A[14]), .B(n31), .CI(n89), .CO(n90), .S(DIFF[14]) );
  inv0d1 U106 ( .I(B[14]), .ZN(n31) );
  ad01d0 U107 ( .A(A[13]), .B(n30), .CI(n88), .CO(n89), .S(DIFF[13]) );
  inv0d1 U108 ( .I(B[13]), .ZN(n30) );
  nr02d0 U109 ( .A1(n21), .A2(A[4]), .ZN(n58) );
  ad01d0 U110 ( .A(A[12]), .B(n29), .CI(n87), .CO(n88), .S(DIFF[12]) );
  inv0d1 U111 ( .I(B[12]), .ZN(n29) );
  ad01d0 U112 ( .A(A[11]), .B(n28), .CI(n86), .CO(n87), .S(DIFF[11]) );
  inv0d1 U113 ( .I(B[11]), .ZN(n28) );
  ad01d0 U114 ( .A(A[10]), .B(n27), .CI(n140), .CO(n86), .S(DIFF[10]) );
  inv0d1 U115 ( .I(B[10]), .ZN(n27) );
  inv0d1 U116 ( .I(n76), .ZN(n77) );
  inv0d1 U117 ( .I(B[9]), .ZN(n26) );
  inv0d1 U118 ( .I(n79), .ZN(n40) );
  inv0d1 U119 ( .I(B[8]), .ZN(n25) );
  nr02d0 U120 ( .A1(n19), .A2(A[2]), .ZN(n49) );
  inv0d1 U121 ( .I(B[2]), .ZN(n19) );
  inv0d1 U122 ( .I(n82), .ZN(n41) );
  inv0d1 U123 ( .I(B[1]), .ZN(n18) );
  nr02d0 U124 ( .A1(n23), .A2(A[6]), .ZN(n68) );
  inv0d1 U125 ( .I(B[6]), .ZN(n23) );
  aoi21d1 U126 ( .B1(n56), .B2(n36), .A(n59), .ZN(n61) );
  aoi21d1 U127 ( .B1(n56), .B2(n65), .A(n64), .ZN(n66) );
  inv0d1 U128 ( .I(n55), .ZN(n56) );
  aoi21d1 U129 ( .B1(n46), .B2(n54), .A(n53), .ZN(n55) );
  inv0d1 U130 ( .I(n46), .ZN(n47) );
  inv0d1 U131 ( .I(B[0]), .ZN(n17) );
  inv0d1 U132 ( .I(n57), .ZN(n59) );
  inv0d1 U133 ( .I(n71), .ZN(n39) );
  inv0d1 U134 ( .I(n52), .ZN(n35) );
  inv0d1 U135 ( .I(n63), .ZN(n37) );
  inv0d1 U136 ( .I(n58), .ZN(n36) );
  inv0d1 U137 ( .I(n49), .ZN(n34) );
  inv0d1 U138 ( .I(B[4]), .ZN(n21) );
  inv0d1 U139 ( .I(n68), .ZN(n38) );
  nr02d0 U140 ( .A1(n63), .A2(n58), .ZN(n65) );
  inv0d1 U141 ( .I(n45), .ZN(n33) );
  inv0d1 U142 ( .I(B[3]), .ZN(n20) );
  aoi21d1 U143 ( .B1(n64), .B2(n73), .A(n72), .ZN(n74) );
  inv0d1 U144 ( .I(B[5]), .ZN(n22) );
  inv0d1 U145 ( .I(B[7]), .ZN(n24) );
endmodule


module BLENDER_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n140;

  nr02d0 U17 ( .A1(n17), .A2(A[0]), .ZN(n43) );
  xn02d1 U18 ( .A1(n17), .A2(A[0]), .ZN(DIFF[0]) );
  nd02d1 U19 ( .A1(n18), .A2(A[1]), .ZN(n44) );
  nd02d1 U22 ( .A1(n33), .A2(n44), .ZN(n91) );
  oai21d1 U23 ( .B1(n45), .B2(n43), .A(n44), .ZN(n46) );
  xr02d1 U25 ( .A1(n91), .A2(n43), .Z(DIFF[1]) );
  nd02d1 U26 ( .A1(n19), .A2(A[2]), .ZN(n48) );
  nr02d0 U27 ( .A1(n19), .A2(A[2]), .ZN(n49) );
  nd02d1 U29 ( .A1(n34), .A2(n48), .ZN(n92) );
  oai21d1 U30 ( .B1(n47), .B2(n49), .A(n48), .ZN(n50) );
  xr02d1 U31 ( .A1(n47), .A2(n92), .Z(DIFF[2]) );
  nd02d1 U32 ( .A1(n20), .A2(A[3]), .ZN(n51) );
  nr02d0 U33 ( .A1(n20), .A2(A[3]), .ZN(n52) );
  nd02d1 U35 ( .A1(n35), .A2(n51), .ZN(n93) );
  oai21d1 U36 ( .B1(n52), .B2(n48), .A(n51), .ZN(n53) );
  nr02d0 U37 ( .A1(n49), .A2(n52), .ZN(n54) );
  xn02d1 U40 ( .A1(n50), .A2(n93), .ZN(DIFF[3]) );
  nd02d1 U41 ( .A1(n21), .A2(A[4]), .ZN(n57) );
  nd02d1 U44 ( .A1(n36), .A2(n57), .ZN(n94) );
  xn02d1 U48 ( .A1(n56), .A2(n94), .ZN(DIFF[4]) );
  nd02d1 U49 ( .A1(n22), .A2(A[5]), .ZN(n62) );
  nd02d1 U52 ( .A1(n37), .A2(n62), .ZN(n95) );
  oai21d1 U53 ( .B1(n63), .B2(n57), .A(n62), .ZN(n64) );
  nr02d0 U54 ( .A1(n58), .A2(n63), .ZN(n65) );
  xr02d1 U56 ( .A1(n61), .A2(n95), .Z(DIFF[5]) );
  nd02d1 U57 ( .A1(n23), .A2(A[6]), .ZN(n67) );
  nd02d1 U60 ( .A1(n38), .A2(n67), .ZN(n96) );
  oai21d1 U61 ( .B1(n66), .B2(n68), .A(n67), .ZN(n69) );
  xr02d1 U62 ( .A1(n66), .A2(n96), .Z(DIFF[6]) );
  nd02d1 U63 ( .A1(n24), .A2(A[7]), .ZN(n70) );
  nd02d1 U66 ( .A1(n39), .A2(n70), .ZN(n97) );
  oai21d1 U67 ( .B1(n71), .B2(n67), .A(n70), .ZN(n72) );
  nr02d0 U68 ( .A1(n71), .A2(n68), .ZN(n73) );
  nd02d1 U70 ( .A1(n65), .A2(n73), .ZN(n75) );
  oai21d1 U71 ( .B1(n55), .B2(n75), .A(n74), .ZN(n76) );
  xn02d1 U73 ( .A1(n69), .A2(n97), .ZN(DIFF[7]) );
  nd02d1 U74 ( .A1(n25), .A2(A[8]), .ZN(n78) );
  nr02d0 U75 ( .A1(n25), .A2(A[8]), .ZN(n79) );
  nd02d1 U77 ( .A1(n40), .A2(n78), .ZN(n98) );
  oai21d1 U78 ( .B1(n77), .B2(n79), .A(n78), .ZN(n80) );
  xr02d1 U79 ( .A1(n77), .A2(n98), .Z(DIFF[8]) );
  nd02d1 U80 ( .A1(n26), .A2(A[9]), .ZN(n81) );
  nr02d0 U81 ( .A1(n26), .A2(A[9]), .ZN(n82) );
  nd02d1 U83 ( .A1(n41), .A2(n81), .ZN(n99) );
  oai21d1 U84 ( .B1(n82), .B2(n78), .A(n81), .ZN(n83) );
  nr02d0 U85 ( .A1(n79), .A2(n82), .ZN(n84) );
  xn02d1 U87 ( .A1(n80), .A2(n99), .ZN(DIFF[9]) );
  xr02d1 U99 ( .A1(n90), .A2(n100), .Z(DIFF[15]) );
  xn02d1 U100 ( .A1(B[15]), .A2(A[15]), .ZN(n100) );
  aor21d1 U101 ( .B1(n76), .B2(n84), .A(n83), .Z(n140) );
  ad01d0 U102 ( .A(A[14]), .B(n31), .CI(n89), .CO(n90), .S(DIFF[14]) );
  inv0d1 U103 ( .I(B[14]), .ZN(n31) );
  ad01d0 U104 ( .A(A[13]), .B(n30), .CI(n88), .CO(n89), .S(DIFF[13]) );
  inv0d1 U105 ( .I(B[13]), .ZN(n30) );
  ad01d0 U106 ( .A(A[12]), .B(n29), .CI(n87), .CO(n88), .S(DIFF[12]) );
  inv0d1 U107 ( .I(B[12]), .ZN(n29) );
  ad01d0 U108 ( .A(A[11]), .B(n28), .CI(n86), .CO(n87), .S(DIFF[11]) );
  inv0d1 U109 ( .I(B[11]), .ZN(n28) );
  ad01d0 U110 ( .A(A[10]), .B(n27), .CI(n140), .CO(n86), .S(DIFF[10]) );
  inv0d1 U111 ( .I(B[10]), .ZN(n27) );
  inv0d1 U112 ( .I(n76), .ZN(n77) );
  inv0d1 U113 ( .I(B[8]), .ZN(n25) );
  inv0d1 U114 ( .I(n79), .ZN(n40) );
  inv0d1 U115 ( .I(n82), .ZN(n41) );
  inv0d1 U116 ( .I(B[2]), .ZN(n19) );
  inv0d1 U117 ( .I(B[9]), .ZN(n26) );
  inv0d1 U118 ( .I(B[3]), .ZN(n20) );
  nr02d0 U119 ( .A1(n21), .A2(A[4]), .ZN(n58) );
  inv0d1 U120 ( .I(B[4]), .ZN(n21) );
  nr02d0 U121 ( .A1(n23), .A2(A[6]), .ZN(n68) );
  inv0d1 U122 ( .I(B[6]), .ZN(n23) );
  inv0d1 U123 ( .I(B[0]), .ZN(n17) );
  nr02d0 U124 ( .A1(n24), .A2(A[7]), .ZN(n71) );
  inv0d1 U125 ( .I(B[7]), .ZN(n24) );
  nr02d0 U126 ( .A1(n18), .A2(A[1]), .ZN(n45) );
  inv0d1 U127 ( .I(B[1]), .ZN(n18) );
  nr02d0 U128 ( .A1(n22), .A2(A[5]), .ZN(n63) );
  inv0d1 U129 ( .I(B[5]), .ZN(n22) );
  inv0d1 U130 ( .I(n57), .ZN(n59) );
  inv0d1 U131 ( .I(n71), .ZN(n39) );
  inv0d1 U132 ( .I(n58), .ZN(n36) );
  inv0d1 U133 ( .I(n68), .ZN(n38) );
  inv0d1 U134 ( .I(n45), .ZN(n33) );
  aoi21d1 U135 ( .B1(n56), .B2(n36), .A(n59), .ZN(n61) );
  aoi21d1 U136 ( .B1(n56), .B2(n65), .A(n64), .ZN(n66) );
  inv0d1 U137 ( .I(n55), .ZN(n56) );
  inv0d1 U138 ( .I(n46), .ZN(n47) );
  aoi21d1 U139 ( .B1(n46), .B2(n54), .A(n53), .ZN(n55) );
  inv0d1 U140 ( .I(n63), .ZN(n37) );
  inv0d1 U141 ( .I(n49), .ZN(n34) );
  inv0d1 U142 ( .I(n52), .ZN(n35) );
  aoi21d1 U143 ( .B1(n64), .B2(n73), .A(n72), .ZN(n74) );
endmodule


module BLENDER_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n128, n129;

  nd02d1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n28) );
  nd02d1 U6 ( .A1(B[1]), .A2(A[1]), .ZN(n30) );
  nd02d1 U9 ( .A1(n18), .A2(n30), .ZN(n78) );
  oai21d1 U10 ( .B1(n31), .B2(n28), .A(n30), .ZN(n32) );
  xr02d1 U12 ( .A1(n78), .A2(n28), .Z(SUM[1]) );
  nd02d1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n34) );
  nr02d0 U14 ( .A1(B[2]), .A2(A[2]), .ZN(n35) );
  nd02d1 U16 ( .A1(n19), .A2(n34), .ZN(n79) );
  oai21d1 U17 ( .B1(n33), .B2(n35), .A(n34), .ZN(n36) );
  xr02d1 U18 ( .A1(n33), .A2(n79), .Z(SUM[2]) );
  nd02d1 U19 ( .A1(B[3]), .A2(A[3]), .ZN(n37) );
  nr02d0 U20 ( .A1(B[3]), .A2(A[3]), .ZN(n38) );
  nd02d1 U22 ( .A1(n20), .A2(n37), .ZN(n80) );
  oai21d1 U23 ( .B1(n38), .B2(n34), .A(n37), .ZN(n39) );
  nr02d0 U24 ( .A1(n35), .A2(n38), .ZN(n40) );
  xn02d1 U27 ( .A1(n36), .A2(n80), .ZN(SUM[3]) );
  nd02d1 U28 ( .A1(B[4]), .A2(A[4]), .ZN(n43) );
  nd02d1 U31 ( .A1(n21), .A2(n43), .ZN(n81) );
  xn02d1 U35 ( .A1(n42), .A2(n81), .ZN(SUM[4]) );
  nd02d1 U36 ( .A1(B[5]), .A2(A[5]), .ZN(n48) );
  nd02d1 U39 ( .A1(n22), .A2(n48), .ZN(n82) );
  oai21d1 U40 ( .B1(n49), .B2(n43), .A(n48), .ZN(n50) );
  xr02d1 U43 ( .A1(n47), .A2(n82), .Z(SUM[5]) );
  nd02d1 U44 ( .A1(B[6]), .A2(A[6]), .ZN(n53) );
  nd02d1 U47 ( .A1(n23), .A2(n53), .ZN(n83) );
  oai21d1 U48 ( .B1(n52), .B2(n54), .A(n53), .ZN(n55) );
  xr02d1 U49 ( .A1(n52), .A2(n83), .Z(SUM[6]) );
  nd02d1 U50 ( .A1(B[7]), .A2(A[7]), .ZN(n56) );
  nr02d0 U51 ( .A1(B[7]), .A2(A[7]), .ZN(n57) );
  nd02d1 U53 ( .A1(n24), .A2(n56), .ZN(n84) );
  oai21d1 U54 ( .B1(n57), .B2(n53), .A(n56), .ZN(n58) );
  nr02d0 U55 ( .A1(n54), .A2(n57), .ZN(n59) );
  nd02d1 U57 ( .A1(n51), .A2(n59), .ZN(n61) );
  oai21d1 U58 ( .B1(n41), .B2(n61), .A(n60), .ZN(n62) );
  xn02d1 U60 ( .A1(n55), .A2(n84), .ZN(SUM[7]) );
  nd02d1 U61 ( .A1(B[8]), .A2(A[8]), .ZN(n64) );
  nr02d0 U62 ( .A1(B[8]), .A2(A[8]), .ZN(n65) );
  nd02d1 U64 ( .A1(n25), .A2(n64), .ZN(n85) );
  oai21d1 U65 ( .B1(n63), .B2(n65), .A(n64), .ZN(n66) );
  xr02d1 U66 ( .A1(n63), .A2(n85), .Z(SUM[8]) );
  nd02d1 U67 ( .A1(B[9]), .A2(A[9]), .ZN(n67) );
  nr02d0 U68 ( .A1(B[9]), .A2(A[9]), .ZN(n68) );
  nd02d1 U70 ( .A1(n26), .A2(n67), .ZN(n86) );
  oai21d1 U71 ( .B1(n68), .B2(n64), .A(n67), .ZN(n69) );
  nr02d0 U72 ( .A1(n65), .A2(n68), .ZN(n70) );
  xn02d1 U74 ( .A1(n66), .A2(n86), .ZN(SUM[9]) );
  xr02d1 U81 ( .A1(B[15]), .A2(A[15]), .Z(n87) );
  ad01d0 U86 ( .A(A[10]), .B(B[10]), .CI(n129), .CO(n72), .S(SUM[10]) );
  an02d1 U87 ( .A1(n128), .A2(n28), .Z(SUM[0]) );
  or02d1 U88 ( .A1(B[0]), .A2(A[0]), .Z(n128) );
  xr02d1 U89 ( .A1(n76), .A2(n87), .Z(SUM[15]) );
  aor21d1 U90 ( .B1(n62), .B2(n70), .A(n69), .Z(n129) );
  ad01d0 U91 ( .A(A[11]), .B(B[11]), .CI(n72), .CO(n73), .S(SUM[11]) );
  ad01d0 U92 ( .A(A[12]), .B(B[12]), .CI(n73), .CO(n74), .S(SUM[12]) );
  ad01d0 U93 ( .A(A[13]), .B(B[13]), .CI(n74), .CO(n75), .S(SUM[13]) );
  ad01d0 U94 ( .A(A[14]), .B(B[14]), .CI(n75), .CO(n76), .S(SUM[14]) );
  nr02d0 U95 ( .A1(B[6]), .A2(A[6]), .ZN(n54) );
  nr02d0 U96 ( .A1(B[5]), .A2(A[5]), .ZN(n49) );
  nr02d0 U97 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  nr02d0 U98 ( .A1(B[4]), .A2(A[4]), .ZN(n44) );
  inv0d1 U99 ( .I(n62), .ZN(n63) );
  inv0d1 U100 ( .I(n65), .ZN(n25) );
  inv0d1 U101 ( .I(n68), .ZN(n26) );
  aoi21d1 U102 ( .B1(n42), .B2(n21), .A(n45), .ZN(n47) );
  aoi21d1 U103 ( .B1(n42), .B2(n51), .A(n50), .ZN(n52) );
  inv0d1 U104 ( .I(n41), .ZN(n42) );
  inv0d1 U105 ( .I(n32), .ZN(n33) );
  aoi21d1 U106 ( .B1(n32), .B2(n40), .A(n39), .ZN(n41) );
  inv0d1 U107 ( .I(n43), .ZN(n45) );
  inv0d1 U108 ( .I(n54), .ZN(n23) );
  inv0d1 U109 ( .I(n31), .ZN(n18) );
  inv0d1 U110 ( .I(n49), .ZN(n22) );
  inv0d1 U111 ( .I(n44), .ZN(n21) );
  inv0d1 U112 ( .I(n35), .ZN(n19) );
  nr02d0 U113 ( .A1(n49), .A2(n44), .ZN(n51) );
  inv0d1 U114 ( .I(n38), .ZN(n20) );
  aoi21d1 U115 ( .B1(n50), .B2(n59), .A(n58), .ZN(n60) );
  inv0d1 U116 ( .I(n57), .ZN(n24) );
endmodule


module BLENDER_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n128, n129;

  nd02d1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n28) );
  nd02d1 U6 ( .A1(B[1]), .A2(A[1]), .ZN(n30) );
  nd02d1 U9 ( .A1(n18), .A2(n30), .ZN(n78) );
  oai21d1 U10 ( .B1(n31), .B2(n28), .A(n30), .ZN(n32) );
  xr02d1 U12 ( .A1(n78), .A2(n28), .Z(SUM[1]) );
  nd02d1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n34) );
  nr02d0 U14 ( .A1(B[2]), .A2(A[2]), .ZN(n35) );
  nd02d1 U16 ( .A1(n19), .A2(n34), .ZN(n79) );
  oai21d1 U17 ( .B1(n33), .B2(n35), .A(n34), .ZN(n36) );
  xr02d1 U18 ( .A1(n33), .A2(n79), .Z(SUM[2]) );
  nd02d1 U19 ( .A1(B[3]), .A2(A[3]), .ZN(n37) );
  nr02d0 U20 ( .A1(B[3]), .A2(A[3]), .ZN(n38) );
  nd02d1 U22 ( .A1(n20), .A2(n37), .ZN(n80) );
  oai21d1 U23 ( .B1(n38), .B2(n34), .A(n37), .ZN(n39) );
  nr02d0 U24 ( .A1(n35), .A2(n38), .ZN(n40) );
  xn02d1 U27 ( .A1(n36), .A2(n80), .ZN(SUM[3]) );
  nd02d1 U28 ( .A1(B[4]), .A2(A[4]), .ZN(n43) );
  nd02d1 U31 ( .A1(n21), .A2(n43), .ZN(n81) );
  xn02d1 U35 ( .A1(n42), .A2(n81), .ZN(SUM[4]) );
  nd02d1 U36 ( .A1(B[5]), .A2(A[5]), .ZN(n48) );
  nd02d1 U39 ( .A1(n22), .A2(n48), .ZN(n82) );
  oai21d1 U40 ( .B1(n49), .B2(n43), .A(n48), .ZN(n50) );
  nr02d0 U41 ( .A1(n44), .A2(n49), .ZN(n51) );
  xr02d1 U43 ( .A1(n47), .A2(n82), .Z(SUM[5]) );
  nd02d1 U44 ( .A1(B[6]), .A2(A[6]), .ZN(n53) );
  nd02d1 U47 ( .A1(n23), .A2(n53), .ZN(n83) );
  oai21d1 U48 ( .B1(n52), .B2(n54), .A(n53), .ZN(n55) );
  xr02d1 U49 ( .A1(n52), .A2(n83), .Z(SUM[6]) );
  nd02d1 U50 ( .A1(B[7]), .A2(A[7]), .ZN(n56) );
  nr02d0 U51 ( .A1(B[7]), .A2(A[7]), .ZN(n57) );
  nd02d1 U53 ( .A1(n24), .A2(n56), .ZN(n84) );
  oai21d1 U54 ( .B1(n57), .B2(n53), .A(n56), .ZN(n58) );
  nr02d0 U55 ( .A1(n54), .A2(n57), .ZN(n59) );
  nd02d1 U57 ( .A1(n51), .A2(n59), .ZN(n61) );
  oai21d1 U58 ( .B1(n41), .B2(n61), .A(n60), .ZN(n62) );
  xn02d1 U60 ( .A1(n55), .A2(n84), .ZN(SUM[7]) );
  nd02d1 U61 ( .A1(B[8]), .A2(A[8]), .ZN(n64) );
  nr02d0 U62 ( .A1(B[8]), .A2(A[8]), .ZN(n65) );
  nd02d1 U64 ( .A1(n25), .A2(n64), .ZN(n85) );
  oai21d1 U65 ( .B1(n63), .B2(n65), .A(n64), .ZN(n66) );
  xr02d1 U66 ( .A1(n63), .A2(n85), .Z(SUM[8]) );
  nd02d1 U67 ( .A1(B[9]), .A2(A[9]), .ZN(n67) );
  nr02d0 U68 ( .A1(B[9]), .A2(A[9]), .ZN(n68) );
  nd02d1 U70 ( .A1(n26), .A2(n67), .ZN(n86) );
  oai21d1 U71 ( .B1(n68), .B2(n64), .A(n67), .ZN(n69) );
  nr02d0 U72 ( .A1(n65), .A2(n68), .ZN(n70) );
  xn02d1 U74 ( .A1(n66), .A2(n86), .ZN(SUM[9]) );
  xr02d1 U81 ( .A1(B[15]), .A2(A[15]), .Z(n87) );
  ad01d0 U86 ( .A(A[10]), .B(B[10]), .CI(n129), .CO(n72), .S(SUM[10]) );
  an02d1 U87 ( .A1(n128), .A2(n28), .Z(SUM[0]) );
  or02d1 U88 ( .A1(B[0]), .A2(A[0]), .Z(n128) );
  xr02d1 U89 ( .A1(n76), .A2(n87), .Z(SUM[15]) );
  aor21d1 U90 ( .B1(n62), .B2(n70), .A(n69), .Z(n129) );
  ad01d0 U91 ( .A(A[13]), .B(B[13]), .CI(n74), .CO(n75), .S(SUM[13]) );
  ad01d0 U92 ( .A(A[11]), .B(B[11]), .CI(n72), .CO(n73), .S(SUM[11]) );
  ad01d0 U93 ( .A(A[12]), .B(B[12]), .CI(n73), .CO(n74), .S(SUM[12]) );
  ad01d0 U94 ( .A(A[14]), .B(B[14]), .CI(n75), .CO(n76), .S(SUM[14]) );
  nr02d0 U95 ( .A1(B[5]), .A2(A[5]), .ZN(n49) );
  nr02d0 U96 ( .A1(B[6]), .A2(A[6]), .ZN(n54) );
  nr02d0 U97 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  nr02d0 U98 ( .A1(B[4]), .A2(A[4]), .ZN(n44) );
  inv0d1 U99 ( .I(n62), .ZN(n63) );
  inv0d1 U100 ( .I(n65), .ZN(n25) );
  inv0d1 U101 ( .I(n68), .ZN(n26) );
  aoi21d1 U102 ( .B1(n42), .B2(n21), .A(n45), .ZN(n47) );
  aoi21d1 U103 ( .B1(n42), .B2(n51), .A(n50), .ZN(n52) );
  inv0d1 U104 ( .I(n41), .ZN(n42) );
  inv0d1 U105 ( .I(n32), .ZN(n33) );
  aoi21d1 U106 ( .B1(n32), .B2(n40), .A(n39), .ZN(n41) );
  inv0d1 U107 ( .I(n43), .ZN(n45) );
  inv0d1 U108 ( .I(n54), .ZN(n23) );
  inv0d1 U109 ( .I(n44), .ZN(n21) );
  inv0d1 U110 ( .I(n31), .ZN(n18) );
  inv0d1 U111 ( .I(n49), .ZN(n22) );
  inv0d1 U112 ( .I(n35), .ZN(n19) );
  inv0d1 U113 ( .I(n38), .ZN(n20) );
  aoi21d1 U114 ( .B1(n50), .B2(n59), .A(n58), .ZN(n60) );
  inv0d1 U115 ( .I(n57), .ZN(n24) );
endmodule


module BLENDER_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n35, n38, n41, n42, n43, n44, n47, n48, n51, n52, n55, n58, n59, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n85, n158;

  or02d1 U3 ( .A1(A[0]), .A2(A[1]), .Z(n35) );
  xn02d1 U4 ( .A1(A[0]), .A2(A[1]), .ZN(SUM[1]) );
  nr02d0 U8 ( .A1(n35), .A2(A[2]), .ZN(n38) );
  xn02d1 U9 ( .A1(n35), .A2(A[2]), .ZN(SUM[2]) );
  nd02d1 U12 ( .A1(A[3]), .A2(A[2]), .ZN(n41) );
  oai21d1 U15 ( .B1(n85), .B2(n42), .A(n41), .ZN(n43) );
  xr02d1 U17 ( .A1(n38), .A2(n42), .Z(SUM[3]) );
  nr02d0 U21 ( .A1(n44), .A2(n47), .ZN(n48) );
  xr02d1 U22 ( .A1(n44), .A2(n47), .Z(SUM[4]) );
  nd02d1 U25 ( .A1(A[4]), .A2(A[5]), .ZN(n51) );
  nr02d0 U26 ( .A1(n44), .A2(n51), .ZN(n52) );
  nd02d1 U30 ( .A1(n52), .A2(A[6]), .ZN(n55) );
  nd02d1 U34 ( .A1(A[6]), .A2(A[7]), .ZN(n58) );
  nr02d0 U35 ( .A1(n51), .A2(n58), .ZN(n59) );
  ah01d0 U39 ( .A(A[8]), .B(n158), .CO(n61), .S(SUM[8]) );
  ah01d0 U40 ( .A(A[9]), .B(n61), .CO(n62), .S(SUM[9]) );
  ah01d0 U41 ( .A(A[10]), .B(n62), .CO(n63), .S(SUM[10]) );
  ah01d0 U42 ( .A(A[11]), .B(n63), .CO(n64), .S(SUM[11]) );
  ah01d0 U43 ( .A(A[12]), .B(n64), .CO(n65), .S(SUM[12]) );
  ah01d0 U44 ( .A(A[13]), .B(n65), .CO(n66), .S(SUM[13]) );
  ah01d0 U45 ( .A(A[14]), .B(n66), .CO(n67), .S(SUM[14]) );
  ah01d0 U46 ( .A(A[15]), .B(n67), .CO(n68), .S(SUM[15]) );
  ah01d0 U47 ( .A(A[16]), .B(n68), .CO(n69), .S(SUM[16]) );
  ah01d0 U48 ( .A(A[17]), .B(n69), .CO(n70), .S(SUM[17]) );
  ah01d0 U49 ( .A(A[18]), .B(n70), .CO(n71), .S(SUM[18]) );
  ah01d0 U50 ( .A(A[19]), .B(n71), .CO(n72), .S(SUM[19]) );
  ah01d0 U51 ( .A(A[20]), .B(n72), .CO(n73), .S(SUM[20]) );
  ah01d0 U52 ( .A(A[21]), .B(n73), .CO(n74), .S(SUM[21]) );
  ah01d0 U53 ( .A(A[22]), .B(n74), .CO(n75), .S(SUM[22]) );
  ah01d0 U54 ( .A(A[23]), .B(n75), .CO(n76), .S(SUM[23]) );
  ah01d0 U55 ( .A(A[24]), .B(n76), .CO(n77), .S(SUM[24]) );
  ah01d0 U56 ( .A(A[25]), .B(n77), .CO(n78), .S(SUM[25]) );
  ah01d0 U57 ( .A(A[26]), .B(n78), .CO(n79), .S(SUM[26]) );
  ah01d0 U58 ( .A(A[27]), .B(n79), .CO(n80), .S(SUM[27]) );
  ah01d0 U59 ( .A(A[28]), .B(n80), .CO(n81), .S(SUM[28]) );
  ah01d0 U60 ( .A(A[29]), .B(n81), .CO(n82), .S(SUM[29]) );
  ah01d0 U61 ( .A(A[30]), .B(n82), .CO(n83), .S(SUM[30]) );
  xr02d1 U62 ( .A1(n83), .A2(A[31]), .Z(SUM[31]) );
  inv0d1 U67 ( .I(n43), .ZN(n44) );
  an02d1 U68 ( .A1(n43), .A2(n59), .Z(n158) );
  inv0d1 U69 ( .I(A[3]), .ZN(n42) );
  inv0d1 U70 ( .I(n35), .ZN(n85) );
  xr02d1 U71 ( .A1(n48), .A2(A[5]), .Z(SUM[5]) );
  xr02d1 U72 ( .A1(n52), .A2(A[6]), .Z(SUM[6]) );
  xn02d1 U73 ( .A1(n55), .A2(A[7]), .ZN(SUM[7]) );
  inv0d1 U74 ( .I(A[4]), .ZN(n47) );
  inv0d1 U75 ( .I(A[0]), .ZN(SUM[0]) );
endmodule


module BLENDER_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n35, n38, n39, n40, n41, n42, n46, n49, n50, n51, n54, n57, n58, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n88, n161;

  ah01d0 U3 ( .A(A[1]), .B(A[0]), .CO(n35), .S(DIFF[1]) );
  nd02d1 U6 ( .A1(n35), .A2(A[2]), .ZN(n38) );
  xn02d1 U7 ( .A1(n35), .A2(n40), .ZN(DIFF[2]) );
  oai21d1 U12 ( .B1(n88), .B2(n40), .A(n39), .ZN(n41) );
  xr02d1 U14 ( .A1(n38), .A2(A[3]), .Z(DIFF[3]) );
  nr02d0 U18 ( .A1(n42), .A2(n50), .ZN(n46) );
  xr02d1 U19 ( .A1(n42), .A2(n50), .Z(DIFF[4]) );
  oai21d1 U25 ( .B1(n42), .B2(n50), .A(n49), .ZN(n51) );
  xn02d1 U26 ( .A1(n46), .A2(A[5]), .ZN(DIFF[5]) );
  nr02d0 U30 ( .A1(n51), .A2(A[6]), .ZN(n54) );
  xn02d1 U31 ( .A1(n51), .A2(A[6]), .ZN(DIFF[6]) );
  nr02d0 U35 ( .A1(A[7]), .A2(A[6]), .ZN(n57) );
  nd02d1 U36 ( .A1(n57), .A2(n49), .ZN(n58) );
  xr02d1 U39 ( .A1(n54), .A2(A[7]), .Z(DIFF[7]) );
  or02d1 U41 ( .A1(n161), .A2(A[8]), .Z(n61) );
  xn02d1 U42 ( .A1(n161), .A2(A[8]), .ZN(DIFF[8]) );
  or02d1 U43 ( .A1(n61), .A2(A[9]), .Z(n62) );
  xn02d1 U44 ( .A1(n61), .A2(A[9]), .ZN(DIFF[9]) );
  or02d1 U45 ( .A1(n62), .A2(A[10]), .Z(n63) );
  xn02d1 U46 ( .A1(n62), .A2(A[10]), .ZN(DIFF[10]) );
  or02d1 U47 ( .A1(n63), .A2(A[11]), .Z(n64) );
  xn02d1 U48 ( .A1(n63), .A2(A[11]), .ZN(DIFF[11]) );
  or02d1 U49 ( .A1(n64), .A2(A[12]), .Z(n65) );
  xn02d1 U50 ( .A1(n64), .A2(A[12]), .ZN(DIFF[12]) );
  or02d1 U51 ( .A1(n65), .A2(A[13]), .Z(n66) );
  xn02d1 U52 ( .A1(n65), .A2(A[13]), .ZN(DIFF[13]) );
  or02d1 U53 ( .A1(n66), .A2(A[14]), .Z(n67) );
  xn02d1 U54 ( .A1(n66), .A2(A[14]), .ZN(DIFF[14]) );
  or02d1 U55 ( .A1(n67), .A2(A[15]), .Z(n68) );
  xn02d1 U56 ( .A1(n67), .A2(A[15]), .ZN(DIFF[15]) );
  or02d1 U57 ( .A1(n68), .A2(A[16]), .Z(n69) );
  xn02d1 U58 ( .A1(n68), .A2(A[16]), .ZN(DIFF[16]) );
  or02d1 U59 ( .A1(n69), .A2(A[17]), .Z(n70) );
  xn02d1 U60 ( .A1(n69), .A2(A[17]), .ZN(DIFF[17]) );
  or02d1 U61 ( .A1(n70), .A2(A[18]), .Z(n71) );
  xn02d1 U62 ( .A1(n70), .A2(A[18]), .ZN(DIFF[18]) );
  or02d1 U63 ( .A1(n71), .A2(A[19]), .Z(n72) );
  xn02d1 U64 ( .A1(n71), .A2(A[19]), .ZN(DIFF[19]) );
  or02d1 U65 ( .A1(n72), .A2(A[20]), .Z(n73) );
  xn02d1 U66 ( .A1(n72), .A2(A[20]), .ZN(DIFF[20]) );
  or02d1 U67 ( .A1(n73), .A2(A[21]), .Z(n74) );
  xn02d1 U68 ( .A1(n73), .A2(A[21]), .ZN(DIFF[21]) );
  or02d1 U69 ( .A1(n74), .A2(A[22]), .Z(n75) );
  xn02d1 U70 ( .A1(n74), .A2(A[22]), .ZN(DIFF[22]) );
  or02d1 U71 ( .A1(n75), .A2(A[23]), .Z(n76) );
  xn02d1 U72 ( .A1(n75), .A2(A[23]), .ZN(DIFF[23]) );
  or02d1 U73 ( .A1(n76), .A2(A[24]), .Z(n77) );
  xn02d1 U74 ( .A1(n76), .A2(A[24]), .ZN(DIFF[24]) );
  or02d1 U75 ( .A1(n77), .A2(A[25]), .Z(n78) );
  xn02d1 U76 ( .A1(n77), .A2(A[25]), .ZN(DIFF[25]) );
  or02d1 U77 ( .A1(n78), .A2(A[26]), .Z(n79) );
  xn02d1 U78 ( .A1(n78), .A2(A[26]), .ZN(DIFF[26]) );
  or02d1 U79 ( .A1(n79), .A2(A[27]), .Z(n80) );
  xn02d1 U80 ( .A1(n79), .A2(A[27]), .ZN(DIFF[27]) );
  or02d1 U81 ( .A1(n80), .A2(A[28]), .Z(n81) );
  xn02d1 U82 ( .A1(n80), .A2(A[28]), .ZN(DIFF[28]) );
  or02d1 U83 ( .A1(n81), .A2(A[29]), .Z(n82) );
  xn02d1 U84 ( .A1(n81), .A2(A[29]), .ZN(DIFF[29]) );
  or02d1 U85 ( .A1(n82), .A2(A[30]), .Z(n83) );
  xn02d1 U86 ( .A1(n82), .A2(A[30]), .ZN(DIFF[30]) );
  xn02d1 U87 ( .A1(n83), .A2(A[31]), .ZN(DIFF[31]) );
  inv0d1 U92 ( .I(n41), .ZN(n42) );
  inv0d1 U93 ( .I(A[3]), .ZN(n39) );
  inv0d1 U94 ( .I(n35), .ZN(n88) );
  inv0d1 U95 ( .I(A[2]), .ZN(n40) );
  aor21d1 U96 ( .B1(n41), .B2(A[4]), .A(n58), .Z(n161) );
  inv0d1 U97 ( .I(A[5]), .ZN(n49) );
  inv0d1 U98 ( .I(A[4]), .ZN(n50) );
  inv0d1 U99 ( .I(A[0]), .ZN(DIFF[0]) );
endmodule


module BLENDER_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n35, n38, n39, n40, n41, n42, n45, n46, n49, n50, n51, n54, n57, n58,
         n59, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n86, n159;

  or02d1 U3 ( .A1(A[0]), .A2(A[1]), .Z(n35) );
  xn02d1 U4 ( .A1(A[0]), .A2(A[1]), .ZN(DIFF[1]) );
  nd02d1 U7 ( .A1(n35), .A2(A[2]), .ZN(n38) );
  xn02d1 U8 ( .A1(n35), .A2(n40), .ZN(DIFF[2]) );
  oai21d1 U13 ( .B1(n86), .B2(n40), .A(n39), .ZN(n41) );
  xr02d1 U15 ( .A1(n38), .A2(A[3]), .Z(DIFF[3]) );
  nd02d1 U20 ( .A1(n42), .A2(n45), .ZN(n46) );
  xr02d1 U21 ( .A1(n42), .A2(A[4]), .Z(DIFF[4]) );
  nd02d1 U24 ( .A1(A[5]), .A2(A[4]), .ZN(n49) );
  oai21d1 U26 ( .B1(n42), .B2(n50), .A(n49), .ZN(n51) );
  xn02d1 U27 ( .A1(n46), .A2(n50), .ZN(DIFF[5]) );
  nd02d1 U30 ( .A1(n51), .A2(A[6]), .ZN(n54) );
  nd02d1 U34 ( .A1(A[6]), .A2(A[7]), .ZN(n57) );
  nr02d0 U35 ( .A1(n57), .A2(n49), .ZN(n58) );
  nr02d0 U36 ( .A1(n57), .A2(n50), .ZN(n59) );
  ah01d0 U40 ( .A(A[8]), .B(n159), .CO(n61), .S(DIFF[8]) );
  ah01d0 U41 ( .A(A[9]), .B(n61), .CO(n62), .S(DIFF[9]) );
  or02d1 U42 ( .A1(n62), .A2(A[10]), .Z(n63) );
  xn02d1 U43 ( .A1(n62), .A2(A[10]), .ZN(DIFF[10]) );
  or02d1 U44 ( .A1(n63), .A2(A[11]), .Z(n64) );
  xn02d1 U45 ( .A1(n63), .A2(A[11]), .ZN(DIFF[11]) );
  or02d1 U46 ( .A1(n64), .A2(A[12]), .Z(n65) );
  xn02d1 U47 ( .A1(n64), .A2(A[12]), .ZN(DIFF[12]) );
  or02d1 U48 ( .A1(n65), .A2(A[13]), .Z(n66) );
  xn02d1 U49 ( .A1(n65), .A2(A[13]), .ZN(DIFF[13]) );
  or02d1 U50 ( .A1(n66), .A2(A[14]), .Z(n67) );
  xn02d1 U51 ( .A1(n66), .A2(A[14]), .ZN(DIFF[14]) );
  or02d1 U52 ( .A1(n67), .A2(A[15]), .Z(n68) );
  xn02d1 U53 ( .A1(n67), .A2(A[15]), .ZN(DIFF[15]) );
  or02d1 U54 ( .A1(n68), .A2(A[16]), .Z(n69) );
  xn02d1 U55 ( .A1(n68), .A2(A[16]), .ZN(DIFF[16]) );
  or02d1 U56 ( .A1(n69), .A2(A[17]), .Z(n70) );
  xn02d1 U57 ( .A1(n69), .A2(A[17]), .ZN(DIFF[17]) );
  or02d1 U58 ( .A1(n70), .A2(A[18]), .Z(n71) );
  xn02d1 U59 ( .A1(n70), .A2(A[18]), .ZN(DIFF[18]) );
  or02d1 U60 ( .A1(n71), .A2(A[19]), .Z(n72) );
  xn02d1 U61 ( .A1(n71), .A2(A[19]), .ZN(DIFF[19]) );
  or02d1 U62 ( .A1(n72), .A2(A[20]), .Z(n73) );
  xn02d1 U63 ( .A1(n72), .A2(A[20]), .ZN(DIFF[20]) );
  or02d1 U64 ( .A1(n73), .A2(A[21]), .Z(n74) );
  xn02d1 U65 ( .A1(n73), .A2(A[21]), .ZN(DIFF[21]) );
  or02d1 U66 ( .A1(n74), .A2(A[22]), .Z(n75) );
  xn02d1 U67 ( .A1(n74), .A2(A[22]), .ZN(DIFF[22]) );
  or02d1 U68 ( .A1(n75), .A2(A[23]), .Z(n76) );
  xn02d1 U69 ( .A1(n75), .A2(A[23]), .ZN(DIFF[23]) );
  or02d1 U70 ( .A1(n76), .A2(A[24]), .Z(n77) );
  xn02d1 U71 ( .A1(n76), .A2(A[24]), .ZN(DIFF[24]) );
  or02d1 U72 ( .A1(n77), .A2(A[25]), .Z(n78) );
  xn02d1 U73 ( .A1(n77), .A2(A[25]), .ZN(DIFF[25]) );
  or02d1 U74 ( .A1(n78), .A2(A[26]), .Z(n79) );
  xn02d1 U75 ( .A1(n78), .A2(A[26]), .ZN(DIFF[26]) );
  or02d1 U76 ( .A1(n79), .A2(A[27]), .Z(n80) );
  xn02d1 U77 ( .A1(n79), .A2(A[27]), .ZN(DIFF[27]) );
  or02d1 U78 ( .A1(n80), .A2(A[28]), .Z(n81) );
  xn02d1 U79 ( .A1(n80), .A2(A[28]), .ZN(DIFF[28]) );
  or02d1 U80 ( .A1(n81), .A2(A[29]), .Z(n82) );
  xn02d1 U81 ( .A1(n81), .A2(A[29]), .ZN(DIFF[29]) );
  or02d1 U82 ( .A1(n82), .A2(A[30]), .Z(n83) );
  xn02d1 U83 ( .A1(n82), .A2(A[30]), .ZN(DIFF[30]) );
  xn02d1 U84 ( .A1(n83), .A2(A[31]), .ZN(DIFF[31]) );
  inv0d1 U89 ( .I(n41), .ZN(n42) );
  aor21d1 U90 ( .B1(n41), .B2(n59), .A(n58), .Z(n159) );
  inv0d1 U91 ( .I(A[3]), .ZN(n39) );
  inv0d1 U92 ( .I(n35), .ZN(n86) );
  inv0d1 U93 ( .I(A[2]), .ZN(n40) );
  inv0d1 U94 ( .I(A[5]), .ZN(n50) );
  inv0d1 U95 ( .I(A[4]), .ZN(n45) );
  xr02d1 U96 ( .A1(n51), .A2(A[6]), .Z(DIFF[6]) );
  xn02d1 U97 ( .A1(n54), .A2(A[7]), .ZN(DIFF[7]) );
  inv0d1 U98 ( .I(A[0]), .ZN(DIFF[0]) );
endmodule


module BLENDER_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n34, n37, n38, n39, n40, n41, n45, n48, n49, n50, n51, n52, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n81, n154;

  or02d1 U3 ( .A1(A[1]), .A2(A[2]), .Z(n34) );
  xn02d1 U4 ( .A1(A[1]), .A2(A[2]), .ZN(SUM[2]) );
  nd02d1 U7 ( .A1(n34), .A2(A[3]), .ZN(n37) );
  xn02d1 U8 ( .A1(n34), .A2(n39), .ZN(SUM[3]) );
  oai21d1 U13 ( .B1(n81), .B2(n39), .A(n38), .ZN(n40) );
  xr02d1 U15 ( .A1(n37), .A2(A[4]), .Z(SUM[4]) );
  nr02d0 U19 ( .A1(n41), .A2(n49), .ZN(n45) );
  xr02d1 U20 ( .A1(n41), .A2(n49), .Z(SUM[5]) );
  oai21d1 U26 ( .B1(n41), .B2(n49), .A(n48), .ZN(n50) );
  xn02d1 U27 ( .A1(n45), .A2(A[6]), .ZN(SUM[6]) );
  nd02d1 U30 ( .A1(n48), .A2(n51), .ZN(n52) );
  xn02d1 U33 ( .A1(n50), .A2(A[7]), .ZN(SUM[7]) );
  ah01d0 U35 ( .A(A[8]), .B(n154), .CO(n55), .S(SUM[8]) );
  ah01d0 U36 ( .A(A[9]), .B(n55), .CO(n56), .S(SUM[9]) );
  ah01d0 U37 ( .A(A[10]), .B(n56), .CO(n57), .S(SUM[10]) );
  ah01d0 U38 ( .A(A[11]), .B(n57), .CO(n58), .S(SUM[11]) );
  ah01d0 U39 ( .A(A[12]), .B(n58), .CO(n59), .S(SUM[12]) );
  ah01d0 U40 ( .A(A[13]), .B(n59), .CO(n60), .S(SUM[13]) );
  ah01d0 U41 ( .A(A[14]), .B(n60), .CO(n61), .S(SUM[14]) );
  ah01d0 U42 ( .A(A[15]), .B(n61), .CO(n62), .S(SUM[15]) );
  ah01d0 U43 ( .A(A[16]), .B(n62), .CO(n63), .S(SUM[16]) );
  ah01d0 U44 ( .A(A[17]), .B(n63), .CO(n64), .S(SUM[17]) );
  ah01d0 U45 ( .A(A[18]), .B(n64), .CO(n65), .S(SUM[18]) );
  ah01d0 U46 ( .A(A[19]), .B(n65), .CO(n66), .S(SUM[19]) );
  ah01d0 U47 ( .A(A[20]), .B(n66), .CO(n67), .S(SUM[20]) );
  ah01d0 U48 ( .A(A[21]), .B(n67), .CO(n68), .S(SUM[21]) );
  ah01d0 U49 ( .A(A[22]), .B(n68), .CO(n69), .S(SUM[22]) );
  ah01d0 U50 ( .A(A[23]), .B(n69), .CO(n70), .S(SUM[23]) );
  ah01d0 U51 ( .A(A[24]), .B(n70), .CO(n71), .S(SUM[24]) );
  ah01d0 U52 ( .A(A[25]), .B(n71), .CO(n72), .S(SUM[25]) );
  ah01d0 U53 ( .A(A[26]), .B(n72), .CO(n73), .S(SUM[26]) );
  ah01d0 U54 ( .A(A[27]), .B(n73), .CO(n74), .S(SUM[27]) );
  ah01d0 U55 ( .A(A[28]), .B(n74), .CO(n75), .S(SUM[28]) );
  ah01d0 U56 ( .A(A[29]), .B(n75), .CO(n76), .S(SUM[29]) );
  ah01d0 U57 ( .A(A[30]), .B(n76), .CO(n77), .S(SUM[30]) );
  xr02d1 U58 ( .A1(n77), .A2(A[31]), .Z(SUM[31]) );
  inv0d1 U63 ( .I(n40), .ZN(n41) );
  inv0d1 U64 ( .I(A[4]), .ZN(n38) );
  inv0d1 U65 ( .I(n34), .ZN(n81) );
  aor21d1 U66 ( .B1(n40), .B2(A[5]), .A(n52), .Z(n154) );
  inv0d1 U67 ( .I(A[3]), .ZN(n39) );
  inv0d1 U68 ( .I(A[6]), .ZN(n48) );
  inv0d1 U69 ( .I(A[7]), .ZN(n51) );
  inv0d1 U70 ( .I(A[1]), .ZN(SUM[1]) );
  inv0d1 U71 ( .I(A[5]), .ZN(n49) );
  bufbd1 U72 ( .I(A[0]), .Z(SUM[0]) );
endmodule


module BLENDER_DW_mult_uns_9 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n741, n743, n747, n748, n753, n756, n758, n759, n760, n761, n763,
         n765, n766, n767, n768, n769, n771, n773, n774, n775, n777, n780,
         n782, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n799, n802, n804, n806, n807, n808, n809,
         n812, n813, n814, n815, n817, n819, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n832, n835, n837, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934;

  nr02d0 U33 ( .A1(n48), .A2(n922), .ZN(product[0]) );
  nr02d0 U34 ( .A1(n49), .A2(n32), .ZN(n65) );
  nr02d0 U35 ( .A1(n50), .A2(n922), .ZN(n66) );
  nr02d0 U36 ( .A1(n51), .A2(n922), .ZN(n67) );
  nr02d0 U37 ( .A1(n52), .A2(n32), .ZN(n68) );
  nr02d0 U38 ( .A1(n53), .A2(n32), .ZN(n69) );
  nr02d0 U39 ( .A1(n54), .A2(n32), .ZN(n70) );
  nr02d0 U40 ( .A1(n55), .A2(n32), .ZN(n71) );
  nr02d0 U41 ( .A1(n56), .A2(n922), .ZN(n72) );
  nr02d0 U42 ( .A1(n57), .A2(n922), .ZN(n73) );
  nr02d0 U43 ( .A1(n58), .A2(n32), .ZN(n74) );
  nr02d0 U44 ( .A1(n59), .A2(n32), .ZN(n75) );
  nr02d0 U45 ( .A1(n60), .A2(n922), .ZN(n76) );
  nr02d0 U46 ( .A1(n61), .A2(n922), .ZN(n77) );
  nr02d0 U47 ( .A1(n62), .A2(n922), .ZN(n78) );
  nr02d0 U48 ( .A1(n63), .A2(n32), .ZN(n79) );
  nr02d0 U49 ( .A1(n48), .A2(n33), .ZN(n80) );
  nr02d0 U50 ( .A1(n49), .A2(n33), .ZN(n81) );
  nr02d0 U51 ( .A1(n50), .A2(n33), .ZN(n82) );
  nr02d0 U52 ( .A1(n51), .A2(n33), .ZN(n83) );
  nr02d0 U53 ( .A1(n52), .A2(n33), .ZN(n84) );
  nr02d0 U54 ( .A1(n53), .A2(n33), .ZN(n85) );
  nr02d0 U55 ( .A1(n54), .A2(n33), .ZN(n86) );
  nr02d0 U56 ( .A1(n55), .A2(n33), .ZN(n87) );
  nr02d0 U57 ( .A1(n56), .A2(n33), .ZN(n88) );
  nr02d0 U58 ( .A1(n57), .A2(n33), .ZN(n89) );
  nr02d0 U59 ( .A1(n58), .A2(n33), .ZN(n90) );
  nr02d0 U60 ( .A1(n59), .A2(n33), .ZN(n91) );
  nr02d0 U61 ( .A1(n60), .A2(n33), .ZN(n92) );
  nr02d0 U62 ( .A1(n61), .A2(n33), .ZN(n93) );
  nr02d0 U63 ( .A1(n62), .A2(n33), .ZN(n94) );
  nr02d0 U64 ( .A1(n63), .A2(n33), .ZN(n95) );
  nr02d0 U65 ( .A1(n48), .A2(n917), .ZN(n96) );
  nr02d0 U66 ( .A1(n49), .A2(n917), .ZN(n97) );
  nr02d0 U67 ( .A1(n50), .A2(n917), .ZN(n98) );
  nr02d0 U68 ( .A1(n51), .A2(n917), .ZN(n99) );
  nr02d0 U69 ( .A1(n52), .A2(n917), .ZN(n100) );
  nr02d0 U70 ( .A1(n53), .A2(n34), .ZN(n101) );
  nr02d0 U71 ( .A1(n54), .A2(n34), .ZN(n102) );
  nr02d0 U72 ( .A1(n55), .A2(n917), .ZN(n103) );
  nr02d0 U73 ( .A1(n56), .A2(n34), .ZN(n104) );
  nr02d0 U74 ( .A1(n57), .A2(n34), .ZN(n105) );
  nr02d0 U75 ( .A1(n58), .A2(n34), .ZN(n106) );
  nr02d0 U76 ( .A1(n59), .A2(n34), .ZN(n107) );
  nr02d0 U77 ( .A1(n60), .A2(n34), .ZN(n108) );
  nr02d0 U78 ( .A1(n61), .A2(n34), .ZN(n109) );
  nr02d0 U79 ( .A1(n62), .A2(n917), .ZN(n110) );
  nr02d0 U80 ( .A1(n63), .A2(n917), .ZN(n111) );
  nr02d0 U81 ( .A1(n48), .A2(n35), .ZN(n112) );
  nr02d0 U82 ( .A1(n49), .A2(n35), .ZN(n113) );
  nr02d0 U83 ( .A1(n50), .A2(n35), .ZN(n114) );
  nr02d0 U84 ( .A1(n51), .A2(n35), .ZN(n115) );
  nr02d0 U85 ( .A1(n52), .A2(n35), .ZN(n116) );
  nr02d0 U86 ( .A1(n53), .A2(n35), .ZN(n117) );
  nr02d0 U87 ( .A1(n54), .A2(n35), .ZN(n118) );
  nr02d0 U88 ( .A1(n55), .A2(n35), .ZN(n119) );
  nr02d0 U89 ( .A1(n56), .A2(n35), .ZN(n120) );
  nr02d0 U90 ( .A1(n57), .A2(n35), .ZN(n121) );
  nr02d0 U91 ( .A1(n58), .A2(n35), .ZN(n122) );
  nr02d0 U92 ( .A1(n59), .A2(n35), .ZN(n123) );
  nr02d0 U93 ( .A1(n60), .A2(n35), .ZN(n124) );
  nr02d0 U94 ( .A1(n61), .A2(n35), .ZN(n125) );
  nr02d0 U95 ( .A1(n62), .A2(n35), .ZN(n126) );
  nr02d0 U96 ( .A1(n63), .A2(n35), .ZN(n127) );
  nr02d0 U97 ( .A1(n48), .A2(n36), .ZN(n128) );
  nr02d0 U98 ( .A1(n49), .A2(n36), .ZN(n129) );
  nr02d0 U99 ( .A1(n50), .A2(n36), .ZN(n130) );
  nr02d0 U100 ( .A1(n51), .A2(n36), .ZN(n131) );
  nr02d0 U101 ( .A1(n52), .A2(n36), .ZN(n132) );
  nr02d0 U102 ( .A1(n53), .A2(n36), .ZN(n133) );
  nr02d0 U104 ( .A1(n55), .A2(n36), .ZN(n135) );
  nr02d0 U105 ( .A1(n56), .A2(n36), .ZN(n136) );
  nr02d0 U106 ( .A1(n57), .A2(n36), .ZN(n137) );
  nr02d0 U107 ( .A1(n58), .A2(n36), .ZN(n138) );
  nr02d0 U108 ( .A1(n59), .A2(n36), .ZN(n139) );
  nr02d0 U109 ( .A1(n60), .A2(n36), .ZN(n140) );
  nr02d0 U110 ( .A1(n61), .A2(n36), .ZN(n141) );
  nr02d0 U111 ( .A1(n62), .A2(n36), .ZN(n142) );
  nr02d0 U112 ( .A1(n63), .A2(n36), .ZN(n143) );
  nr02d0 U113 ( .A1(n48), .A2(n37), .ZN(n144) );
  nr02d0 U114 ( .A1(n49), .A2(n913), .ZN(n145) );
  nr02d0 U115 ( .A1(n50), .A2(n37), .ZN(n146) );
  nr02d0 U116 ( .A1(n51), .A2(n37), .ZN(n147) );
  nr02d0 U117 ( .A1(n52), .A2(n37), .ZN(n148) );
  nr02d0 U118 ( .A1(n53), .A2(n37), .ZN(n149) );
  nr02d0 U119 ( .A1(n54), .A2(n37), .ZN(n150) );
  nr02d0 U120 ( .A1(n55), .A2(n37), .ZN(n151) );
  nr02d0 U121 ( .A1(n56), .A2(n37), .ZN(n152) );
  nr02d0 U122 ( .A1(n57), .A2(n913), .ZN(n153) );
  nr02d0 U123 ( .A1(n58), .A2(n913), .ZN(n154) );
  nr02d0 U124 ( .A1(n59), .A2(n913), .ZN(n155) );
  nr02d0 U125 ( .A1(n60), .A2(n913), .ZN(n156) );
  nr02d0 U126 ( .A1(n61), .A2(n913), .ZN(n157) );
  nr02d0 U127 ( .A1(n62), .A2(n913), .ZN(n158) );
  nr02d0 U128 ( .A1(n63), .A2(n913), .ZN(n159) );
  nr02d0 U129 ( .A1(n48), .A2(n38), .ZN(n160) );
  nr02d0 U130 ( .A1(n49), .A2(n38), .ZN(n161) );
  nr02d0 U131 ( .A1(n50), .A2(n38), .ZN(n162) );
  nr02d0 U132 ( .A1(n51), .A2(n38), .ZN(n163) );
  nr02d0 U133 ( .A1(n52), .A2(n38), .ZN(n164) );
  nr02d0 U134 ( .A1(n53), .A2(n38), .ZN(n165) );
  nr02d0 U136 ( .A1(n55), .A2(n38), .ZN(n167) );
  nr02d0 U137 ( .A1(n56), .A2(n916), .ZN(n168) );
  nr02d0 U138 ( .A1(n57), .A2(n916), .ZN(n169) );
  nr02d0 U139 ( .A1(n58), .A2(n916), .ZN(n170) );
  nr02d0 U140 ( .A1(n59), .A2(n916), .ZN(n171) );
  nr02d0 U141 ( .A1(n60), .A2(n916), .ZN(n172) );
  nr02d0 U142 ( .A1(n61), .A2(n916), .ZN(n173) );
  nr02d0 U143 ( .A1(n62), .A2(n916), .ZN(n174) );
  nr02d0 U144 ( .A1(n63), .A2(n916), .ZN(n175) );
  nr02d0 U145 ( .A1(n48), .A2(n39), .ZN(n176) );
  nr02d0 U146 ( .A1(n49), .A2(n39), .ZN(n177) );
  nr02d0 U147 ( .A1(n50), .A2(n39), .ZN(n178) );
  nr02d0 U148 ( .A1(n51), .A2(n39), .ZN(n179) );
  nr02d0 U149 ( .A1(n52), .A2(n39), .ZN(n180) );
  nr02d0 U150 ( .A1(n53), .A2(n39), .ZN(n181) );
  nr02d0 U151 ( .A1(n54), .A2(n39), .ZN(n182) );
  nr02d0 U152 ( .A1(n55), .A2(n39), .ZN(n183) );
  nr02d0 U153 ( .A1(n56), .A2(n39), .ZN(n184) );
  nr02d0 U154 ( .A1(n57), .A2(n39), .ZN(n185) );
  nr02d0 U155 ( .A1(n58), .A2(n39), .ZN(n186) );
  nr02d0 U156 ( .A1(n59), .A2(n39), .ZN(n187) );
  nr02d0 U157 ( .A1(n60), .A2(n39), .ZN(n188) );
  nr02d0 U158 ( .A1(n61), .A2(n39), .ZN(n189) );
  nr02d0 U159 ( .A1(n62), .A2(n39), .ZN(n190) );
  nr02d0 U160 ( .A1(n63), .A2(n39), .ZN(n191) );
  nr02d0 U161 ( .A1(n48), .A2(n40), .ZN(n192) );
  nr02d0 U162 ( .A1(n49), .A2(n40), .ZN(n193) );
  nr02d0 U163 ( .A1(n50), .A2(n40), .ZN(n194) );
  nr02d0 U164 ( .A1(n51), .A2(n40), .ZN(n195) );
  nr02d0 U165 ( .A1(n52), .A2(n40), .ZN(n196) );
  nr02d0 U166 ( .A1(n53), .A2(n40), .ZN(n197) );
  nr02d0 U167 ( .A1(n54), .A2(n40), .ZN(n198) );
  nr02d0 U168 ( .A1(n55), .A2(n40), .ZN(n199) );
  nr02d0 U169 ( .A1(n56), .A2(n40), .ZN(n200) );
  nr02d0 U170 ( .A1(n57), .A2(n40), .ZN(n201) );
  nr02d0 U171 ( .A1(n58), .A2(n40), .ZN(n202) );
  nr02d0 U172 ( .A1(n911), .A2(n40), .ZN(n203) );
  nr02d0 U173 ( .A1(n910), .A2(n40), .ZN(n204) );
  nr02d0 U174 ( .A1(n61), .A2(n40), .ZN(n205) );
  nr02d0 U175 ( .A1(n62), .A2(n40), .ZN(n206) );
  nr02d0 U176 ( .A1(n63), .A2(n40), .ZN(n207) );
  nr02d0 U177 ( .A1(n48), .A2(n41), .ZN(n208) );
  nr02d0 U178 ( .A1(n49), .A2(n41), .ZN(n209) );
  nr02d0 U179 ( .A1(n50), .A2(n41), .ZN(n210) );
  nr02d0 U180 ( .A1(n51), .A2(n41), .ZN(n211) );
  nr02d0 U181 ( .A1(n52), .A2(n41), .ZN(n212) );
  nr02d0 U182 ( .A1(n53), .A2(n41), .ZN(n213) );
  nr02d0 U183 ( .A1(n54), .A2(n41), .ZN(n214) );
  nr02d0 U184 ( .A1(n55), .A2(n41), .ZN(n215) );
  nr02d0 U185 ( .A1(n56), .A2(n915), .ZN(n216) );
  nr02d0 U186 ( .A1(n57), .A2(n915), .ZN(n217) );
  nr02d0 U187 ( .A1(n58), .A2(n915), .ZN(n218) );
  nr02d0 U188 ( .A1(n911), .A2(n915), .ZN(n219) );
  nr02d0 U189 ( .A1(n910), .A2(n915), .ZN(n220) );
  nr02d0 U190 ( .A1(n61), .A2(n915), .ZN(n221) );
  nr02d0 U191 ( .A1(n62), .A2(n915), .ZN(n222) );
  nr02d0 U192 ( .A1(n63), .A2(n915), .ZN(n223) );
  nr02d0 U193 ( .A1(n48), .A2(n42), .ZN(n224) );
  nr02d0 U194 ( .A1(n49), .A2(n42), .ZN(n225) );
  nr02d0 U195 ( .A1(n50), .A2(n42), .ZN(n226) );
  nr02d0 U196 ( .A1(n51), .A2(n42), .ZN(n227) );
  nr02d0 U197 ( .A1(n52), .A2(n42), .ZN(n228) );
  nr02d0 U198 ( .A1(n53), .A2(n42), .ZN(n229) );
  nr02d0 U199 ( .A1(n54), .A2(n42), .ZN(n230) );
  nr02d0 U200 ( .A1(n55), .A2(n42), .ZN(n231) );
  nr02d0 U201 ( .A1(n56), .A2(n912), .ZN(n232) );
  nr02d0 U202 ( .A1(n57), .A2(n912), .ZN(n233) );
  nr02d0 U203 ( .A1(n58), .A2(n912), .ZN(n234) );
  nr02d0 U204 ( .A1(n911), .A2(n912), .ZN(n235) );
  nr02d0 U205 ( .A1(n910), .A2(n912), .ZN(n236) );
  nr02d0 U206 ( .A1(n61), .A2(n912), .ZN(n237) );
  nr02d0 U207 ( .A1(n62), .A2(n912), .ZN(n238) );
  nr02d0 U208 ( .A1(n63), .A2(n912), .ZN(n239) );
  nr02d0 U209 ( .A1(n48), .A2(n43), .ZN(n240) );
  nr02d0 U210 ( .A1(n49), .A2(n43), .ZN(n241) );
  nr02d0 U211 ( .A1(n50), .A2(n43), .ZN(n242) );
  nr02d0 U212 ( .A1(n51), .A2(n43), .ZN(n243) );
  nr02d0 U213 ( .A1(n52), .A2(n43), .ZN(n244) );
  nr02d0 U214 ( .A1(n53), .A2(n43), .ZN(n245) );
  nr02d0 U215 ( .A1(n54), .A2(n43), .ZN(n246) );
  nr02d0 U216 ( .A1(n55), .A2(n43), .ZN(n247) );
  nr02d0 U217 ( .A1(n56), .A2(n43), .ZN(n248) );
  nr02d0 U218 ( .A1(n57), .A2(n43), .ZN(n249) );
  nr02d0 U219 ( .A1(n58), .A2(n43), .ZN(n250) );
  nr02d0 U220 ( .A1(n911), .A2(n43), .ZN(n251) );
  nr02d0 U221 ( .A1(n910), .A2(n43), .ZN(n252) );
  nr02d0 U222 ( .A1(n61), .A2(n43), .ZN(n253) );
  nr02d0 U223 ( .A1(n62), .A2(n43), .ZN(n254) );
  nr02d0 U224 ( .A1(n63), .A2(n43), .ZN(n255) );
  nr02d0 U225 ( .A1(n48), .A2(n44), .ZN(n256) );
  nr02d0 U226 ( .A1(n49), .A2(n44), .ZN(n257) );
  nr02d0 U227 ( .A1(n50), .A2(n44), .ZN(n258) );
  nr02d0 U228 ( .A1(n51), .A2(n44), .ZN(n259) );
  nr02d0 U229 ( .A1(n52), .A2(n44), .ZN(n260) );
  nr02d0 U230 ( .A1(n53), .A2(n44), .ZN(n261) );
  nr02d0 U231 ( .A1(n54), .A2(n44), .ZN(n262) );
  nr02d0 U232 ( .A1(n55), .A2(n44), .ZN(n263) );
  nr02d0 U233 ( .A1(n56), .A2(n44), .ZN(n264) );
  nr02d0 U234 ( .A1(n57), .A2(n44), .ZN(n265) );
  nr02d0 U235 ( .A1(n58), .A2(n44), .ZN(n266) );
  nr02d0 U236 ( .A1(n911), .A2(n44), .ZN(n267) );
  nr02d0 U237 ( .A1(n910), .A2(n44), .ZN(n268) );
  nr02d0 U238 ( .A1(n61), .A2(n44), .ZN(n269) );
  nr02d0 U239 ( .A1(n62), .A2(n44), .ZN(n270) );
  nr02d0 U240 ( .A1(n63), .A2(n44), .ZN(n271) );
  nr02d0 U241 ( .A1(n48), .A2(n45), .ZN(n272) );
  nr02d0 U242 ( .A1(n49), .A2(n45), .ZN(n273) );
  nr02d0 U243 ( .A1(n50), .A2(n45), .ZN(n274) );
  nr02d0 U244 ( .A1(n51), .A2(n45), .ZN(n275) );
  nr02d0 U245 ( .A1(n52), .A2(n45), .ZN(n276) );
  nr02d0 U246 ( .A1(n53), .A2(n45), .ZN(n277) );
  nr02d0 U247 ( .A1(n54), .A2(n45), .ZN(n278) );
  nr02d0 U248 ( .A1(n55), .A2(n45), .ZN(n279) );
  nr02d0 U249 ( .A1(n56), .A2(n914), .ZN(n280) );
  nr02d0 U250 ( .A1(n57), .A2(n914), .ZN(n281) );
  nr02d0 U251 ( .A1(n58), .A2(n914), .ZN(n282) );
  nr02d0 U252 ( .A1(n911), .A2(n914), .ZN(n283) );
  nr02d0 U253 ( .A1(n910), .A2(n914), .ZN(n284) );
  nr02d0 U254 ( .A1(n61), .A2(n914), .ZN(n285) );
  nr02d0 U255 ( .A1(n62), .A2(n914), .ZN(n286) );
  nr02d0 U256 ( .A1(n63), .A2(n914), .ZN(n287) );
  nr02d0 U257 ( .A1(n48), .A2(n46), .ZN(n288) );
  nr02d0 U258 ( .A1(n49), .A2(n46), .ZN(n289) );
  nr02d0 U259 ( .A1(n50), .A2(n46), .ZN(n290) );
  nr02d0 U260 ( .A1(n51), .A2(n46), .ZN(n291) );
  nr02d0 U261 ( .A1(n52), .A2(n46), .ZN(n292) );
  nr02d0 U262 ( .A1(n53), .A2(n46), .ZN(n293) );
  nr02d0 U263 ( .A1(n54), .A2(n46), .ZN(n294) );
  nr02d0 U264 ( .A1(n55), .A2(n46), .ZN(n295) );
  nr02d0 U265 ( .A1(n56), .A2(n46), .ZN(n296) );
  nr02d0 U266 ( .A1(n57), .A2(n46), .ZN(n297) );
  nr02d0 U267 ( .A1(n58), .A2(n46), .ZN(n298) );
  nr02d0 U268 ( .A1(n911), .A2(n46), .ZN(n299) );
  nr02d0 U269 ( .A1(n910), .A2(n46), .ZN(n300) );
  nr02d0 U270 ( .A1(n61), .A2(n46), .ZN(n301) );
  nr02d0 U271 ( .A1(n62), .A2(n46), .ZN(n302) );
  nr02d0 U272 ( .A1(n63), .A2(n46), .ZN(n303) );
  nr02d0 U273 ( .A1(n48), .A2(n47), .ZN(n304) );
  nr02d0 U274 ( .A1(n49), .A2(n47), .ZN(n305) );
  nr02d0 U275 ( .A1(n50), .A2(n47), .ZN(n306) );
  nr02d0 U276 ( .A1(n51), .A2(n47), .ZN(n307) );
  nr02d0 U277 ( .A1(n52), .A2(n47), .ZN(n308) );
  nr02d0 U278 ( .A1(n53), .A2(n47), .ZN(n309) );
  nr02d0 U279 ( .A1(n54), .A2(n47), .ZN(n310) );
  nr02d0 U280 ( .A1(n55), .A2(n47), .ZN(n311) );
  nr02d0 U281 ( .A1(n56), .A2(n47), .ZN(n312) );
  nr02d0 U282 ( .A1(n57), .A2(n47), .ZN(n313) );
  nr02d0 U283 ( .A1(n58), .A2(n47), .ZN(n314) );
  nr02d0 U284 ( .A1(n911), .A2(n47), .ZN(n315) );
  nr02d0 U285 ( .A1(n910), .A2(n47), .ZN(n316) );
  nr02d0 U286 ( .A1(n61), .A2(n47), .ZN(n317) );
  nr02d0 U287 ( .A1(n62), .A2(n47), .ZN(n318) );
  nr02d0 U288 ( .A1(n63), .A2(n47), .ZN(n319) );
  ah01d0 U289 ( .A(n66), .B(n81), .CO(n321), .S(n320) );
  ah01d0 U290 ( .A(n97), .B(n112), .CO(n323), .S(n322) );
  ah01d0 U292 ( .A(n113), .B(n128), .CO(n327), .S(n326) );
  ah01d0 U295 ( .A(n129), .B(n144), .CO(n333), .S(n332) );
  ah01d0 U299 ( .A(n145), .B(n160), .CO(n341), .S(n340) );
  ah01d0 U304 ( .A(n161), .B(n176), .CO(n351), .S(n350) );
  ah01d0 U310 ( .A(n177), .B(n192), .CO(n363), .S(n362) );
  ah01d0 U317 ( .A(n193), .B(n208), .CO(n377), .S(n376) );
  ah01d0 U325 ( .A(n209), .B(n224), .CO(n393), .S(n392) );
  ah01d0 U334 ( .A(n225), .B(n240), .CO(n411), .S(n410) );
  ah01d0 U344 ( .A(n241), .B(n256), .CO(n431), .S(n430) );
  ah01d0 U355 ( .A(n257), .B(n272), .CO(n453), .S(n452) );
  ah01d0 U367 ( .A(n273), .B(n288), .CO(n477), .S(n476) );
  ah01d0 U380 ( .A(n289), .B(n304), .CO(n503), .S(n502) );
  ah01d0 U394 ( .A(n290), .B(n305), .CO(n531), .S(n530) );
  nd02d1 U499 ( .A1(n65), .A2(n80), .ZN(n756) );
  nd02d1 U504 ( .A1(n320), .A2(n96), .ZN(n758) );
  nr02d0 U505 ( .A1(n320), .A2(n96), .ZN(n759) );
  nd02d1 U507 ( .A1(n741), .A2(n758), .ZN(n857) );
  oai21d1 U508 ( .B1(n759), .B2(n756), .A(n758), .ZN(n760) );
  xr02d1 U509 ( .A1(n857), .A2(n756), .Z(product[2]) );
  nd02d1 U510 ( .A1(n324), .A2(n322), .ZN(n761) );
  nd02d1 U513 ( .A1(n934), .A2(n761), .ZN(n858) );
  xn02d1 U517 ( .A1(n858), .A2(n760), .ZN(product[3]) );
  nd02d1 U518 ( .A1(n330), .A2(n325), .ZN(n766) );
  nr02d0 U519 ( .A1(n330), .A2(n325), .ZN(n767) );
  nd02d1 U521 ( .A1(n743), .A2(n766), .ZN(n859) );
  oai21d1 U522 ( .B1(n767), .B2(n765), .A(n766), .ZN(n768) );
  xr02d1 U523 ( .A1(n859), .A2(n765), .Z(product[4]) );
  nd02d1 U524 ( .A1(n338), .A2(n331), .ZN(n769) );
  nd02d1 U527 ( .A1(n933), .A2(n769), .ZN(n860) );
  xn02d1 U532 ( .A1(n860), .A2(n768), .ZN(product[5]) );
  nd02d1 U533 ( .A1(n348), .A2(n339), .ZN(n775) );
  nd02d1 U536 ( .A1(n931), .A2(n775), .ZN(n861) );
  xn02d1 U540 ( .A1(n861), .A2(n774), .ZN(product[6]) );
  nd02d1 U541 ( .A1(n360), .A2(n349), .ZN(n780) );
  nd02d1 U544 ( .A1(n932), .A2(n780), .ZN(n862) );
  nd02d1 U548 ( .A1(n932), .A2(n931), .ZN(n785) );
  oai21d1 U549 ( .B1(n785), .B2(n773), .A(n784), .ZN(n786) );
  nd02d1 U552 ( .A1(n374), .A2(n361), .ZN(n788) );
  nr02d0 U553 ( .A1(n374), .A2(n361), .ZN(n789) );
  nd02d1 U555 ( .A1(n747), .A2(n788), .ZN(n863) );
  oai21d1 U556 ( .B1(n787), .B2(n789), .A(n788), .ZN(n790) );
  xr02d1 U557 ( .A1(n787), .A2(n863), .Z(product[8]) );
  nd02d1 U558 ( .A1(n390), .A2(n375), .ZN(n791) );
  nr02d0 U559 ( .A1(n390), .A2(n375), .ZN(n792) );
  nd02d1 U561 ( .A1(n748), .A2(n791), .ZN(n864) );
  oai21d1 U562 ( .B1(n792), .B2(n788), .A(n791), .ZN(n793) );
  nr02d0 U563 ( .A1(n792), .A2(n789), .ZN(n794) );
  xn02d1 U566 ( .A1(n790), .A2(n864), .ZN(product[9]) );
  nd02d1 U567 ( .A1(n408), .A2(n391), .ZN(n797) );
  nd02d1 U570 ( .A1(n928), .A2(n797), .ZN(n865) );
  xn02d1 U574 ( .A1(n796), .A2(n865), .ZN(product[10]) );
  nd02d1 U575 ( .A1(n428), .A2(n409), .ZN(n802) );
  nd02d1 U578 ( .A1(n929), .A2(n802), .ZN(n866) );
  nd02d1 U582 ( .A1(n929), .A2(n928), .ZN(n807) );
  oai21d1 U583 ( .B1(n795), .B2(n807), .A(n806), .ZN(n808) );
  nd02d1 U586 ( .A1(n450), .A2(n429), .ZN(n814) );
  nr02d0 U587 ( .A1(n450), .A2(n429), .ZN(n815) );
  xr02d1 U595 ( .A1(n809), .A2(n867), .Z(product[12]) );
  nd02d1 U599 ( .A1(n925), .A2(n817), .ZN(n868) );
  oai21d1 U604 ( .B1(n809), .B2(n822), .A(n821), .ZN(n823) );
  nd02d1 U606 ( .A1(n500), .A2(n475), .ZN(n824) );
  nr02d0 U607 ( .A1(n500), .A2(n475), .ZN(n825) );
  nd02d1 U609 ( .A1(n753), .A2(n824), .ZN(n869) );
  oai21d1 U610 ( .B1(n821), .B2(n825), .A(n824), .ZN(n826) );
  nr02d0 U611 ( .A1(n822), .A2(n825), .ZN(n827) );
  xn02d1 U614 ( .A1(n823), .A2(n869), .ZN(product[14]) );
  nd02d1 U615 ( .A1(n528), .A2(n501), .ZN(n830) );
  nd02d1 U618 ( .A1(n924), .A2(n830), .ZN(n870) );
  xn02d1 U622 ( .A1(n829), .A2(n870), .ZN(product[15]) );
  nd02d1 U623 ( .A1(n556), .A2(n529), .ZN(n835) );
  nd02d1 U626 ( .A1(n926), .A2(n835), .ZN(n871) );
  nd02d1 U630 ( .A1(n926), .A2(n924), .ZN(n840) );
  oai21d1 U631 ( .B1(n828), .B2(n840), .A(n839), .ZN(n841) );
  invbd2 U650 ( .I(a[12]), .ZN(n44) );
  invbd2 U651 ( .I(b[6]), .ZN(n54) );
  invbd2 U652 ( .I(b[2]), .ZN(n50) );
  invbd2 U653 ( .I(b[9]), .ZN(n57) );
  an02d1 U654 ( .A1(n921), .A2(n920), .Z(n908) );
  nd02d1 U655 ( .A1(n474), .A2(n451), .ZN(n817) );
  or02d1 U656 ( .A1(n65), .A2(n80), .Z(n909) );
  ad01d1 U657 ( .A(n736), .B(n733), .CI(n852), .CO(n853), .S(product[28]) );
  inv0d1 U658 ( .I(b[12]), .ZN(n910) );
  ad01d0 U659 ( .A(n719), .B(n726), .CI(n850), .CO(n851), .S(product[26]) );
  ad01d0 U660 ( .A(n732), .B(n727), .CI(n851), .CO(n852), .S(product[27]) );
  inv0d1 U661 ( .I(b[11]), .ZN(n911) );
  inv0d1 U662 ( .I(b[11]), .ZN(n59) );
  inv0d1 U663 ( .I(a[10]), .ZN(n912) );
  inv0d1 U664 ( .I(a[5]), .ZN(n913) );
  inv0d1 U665 ( .I(a[5]), .ZN(n37) );
  inv0d1 U666 ( .I(a[13]), .ZN(n914) );
  inv0d1 U667 ( .I(a[9]), .ZN(n915) );
  inv0d1 U668 ( .I(a[9]), .ZN(n41) );
  inv0d1 U669 ( .I(a[6]), .ZN(n916) );
  nd02d1 U670 ( .A1(n919), .A2(n908), .ZN(n447) );
  inv0d1 U671 ( .I(a[2]), .ZN(n917) );
  nr02d0 U672 ( .A1(n54), .A2(n38), .ZN(n166) );
  nr02d0 U673 ( .A1(n54), .A2(n36), .ZN(n134) );
  inv0d1 U674 ( .I(a[11]), .ZN(n43) );
  inv0d1 U675 ( .I(a[1]), .ZN(n33) );
  inv0d1 U676 ( .I(a[2]), .ZN(n34) );
  inv0d0 U677 ( .I(n828), .ZN(n829) );
  nd02d0 U678 ( .A1(n925), .A2(n813), .ZN(n822) );
  xr02d1 U679 ( .A1(n918), .A2(n868), .Z(product[13]) );
  ora21d1 U680 ( .B1(n809), .B2(n815), .A(n814), .Z(n918) );
  nd02d0 U681 ( .A1(n813), .A2(n814), .ZN(n867) );
  ad01d0 U682 ( .A(n430), .B(n413), .CI(n417), .CO(n441), .S(n440) );
  ad01d0 U683 ( .A(n395), .B(n399), .CI(n397), .CO(n421), .S(n420) );
  ad01d0 U684 ( .A(n416), .B(n412), .CI(n414), .CO(n423), .S(n422) );
  xr03d1 U685 ( .A1(n440), .A2(n421), .A3(n423), .Z(n446) );
  nd02d1 U686 ( .A1(n440), .A2(n423), .ZN(n919) );
  nd02d1 U687 ( .A1(n440), .A2(n421), .ZN(n920) );
  nd02d1 U688 ( .A1(n423), .A2(n421), .ZN(n921) );
  inv0d1 U689 ( .I(a[0]), .ZN(n922) );
  inv0d1 U690 ( .I(n830), .ZN(n832) );
  aoi21d1 U691 ( .B1(n808), .B2(n827), .A(n826), .ZN(n828) );
  inv0d1 U692 ( .I(n835), .ZN(n837) );
  xn02d1 U693 ( .A1(n923), .A2(n871), .ZN(product[16]) );
  aor21d1 U694 ( .B1(n829), .B2(n924), .A(n832), .Z(n923) );
  inv0d1 U695 ( .I(n825), .ZN(n753) );
  inv0d1 U696 ( .I(n808), .ZN(n809) );
  inv0d1 U697 ( .I(n795), .ZN(n796) );
  ad01d0 U698 ( .A(n583), .B(n606), .CI(n842), .CO(n843), .S(product[18]) );
  ad01d0 U699 ( .A(n607), .B(n628), .CI(n843), .CO(n844), .S(product[19]) );
  ad01d0 U700 ( .A(n629), .B(n648), .CI(n844), .CO(n845), .S(product[20]) );
  ad01d0 U701 ( .A(n557), .B(n582), .CI(n841), .CO(n842), .S(product[17]) );
  aoi21d1 U702 ( .B1(n926), .B2(n832), .A(n837), .ZN(n839) );
  aoi21d1 U703 ( .B1(n929), .B2(n799), .A(n804), .ZN(n806) );
  inv0d1 U704 ( .I(n802), .ZN(n804) );
  or02d1 U705 ( .A1(n528), .A2(n501), .Z(n924) );
  or02d1 U706 ( .A1(n474), .A2(n451), .Z(n925) );
  or02d1 U707 ( .A1(n556), .A2(n529), .Z(n926) );
  inv0d1 U708 ( .I(n815), .ZN(n813) );
  inv0d1 U709 ( .I(n797), .ZN(n799) );
  aoi21d1 U710 ( .B1(n786), .B2(n794), .A(n793), .ZN(n795) );
  aoi21d1 U711 ( .B1(n925), .B2(n812), .A(n819), .ZN(n821) );
  inv0d1 U712 ( .I(n814), .ZN(n812) );
  inv0d1 U713 ( .I(n817), .ZN(n819) );
  inv0d1 U714 ( .I(n792), .ZN(n748) );
  inv0d1 U715 ( .I(n789), .ZN(n747) );
  xn02d1 U716 ( .A1(n927), .A2(n866), .ZN(product[11]) );
  aor21d1 U717 ( .B1(n796), .B2(n928), .A(n799), .Z(n927) );
  inv0d1 U718 ( .I(n786), .ZN(n787) );
  inv0d1 U719 ( .I(n773), .ZN(n774) );
  ad01d0 U720 ( .A(n427), .B(n446), .CI(n448), .CO(n451), .S(n450) );
  ad01d0 U721 ( .A(n470), .B(n449), .CI(n472), .CO(n475), .S(n474) );
  ad01d0 U722 ( .A(n524), .B(n499), .CI(n526), .CO(n529), .S(n528) );
  ad01d0 U723 ( .A(n552), .B(n527), .CI(n554), .CO(n557), .S(n556) );
  ad01d0 U724 ( .A(n496), .B(n473), .CI(n498), .CO(n501), .S(n500) );
  ad01d0 U725 ( .A(n649), .B(n666), .CI(n845), .CO(n846), .S(product[21]) );
  ad01d0 U726 ( .A(n667), .B(n682), .CI(n846), .CO(n847), .S(product[22]) );
  ad01d0 U727 ( .A(n683), .B(n696), .CI(n847), .CO(n848), .S(product[23]) );
  ad01d0 U728 ( .A(n697), .B(n708), .CI(n848), .CO(n849), .S(product[24]) );
  ad01d0 U729 ( .A(n709), .B(n718), .CI(n849), .CO(n850), .S(product[25]) );
  aoi21d1 U730 ( .B1(n932), .B2(n777), .A(n782), .ZN(n784) );
  inv0d1 U731 ( .I(n780), .ZN(n782) );
  or02d1 U732 ( .A1(n408), .A2(n391), .Z(n928) );
  or02d1 U733 ( .A1(n428), .A2(n409), .Z(n929) );
  inv0d1 U734 ( .I(n775), .ZN(n777) );
  aoi21d1 U735 ( .B1(n768), .B2(n933), .A(n771), .ZN(n773) );
  inv0d1 U736 ( .I(n769), .ZN(n771) );
  ad01d0 U737 ( .A(n578), .B(n555), .CI(n580), .CO(n583), .S(n582) );
  ad01d0 U738 ( .A(n602), .B(n581), .CI(n604), .CO(n607), .S(n606) );
  ad01d0 U739 ( .A(n624), .B(n605), .CI(n626), .CO(n629), .S(n628) );
  ad01d0 U740 ( .A(n551), .B(n576), .CI(n553), .CO(n581), .S(n580) );
  ad01d0 U741 ( .A(n577), .B(n600), .CI(n579), .CO(n605), .S(n604) );
  ad01d0 U742 ( .A(n601), .B(n622), .CI(n603), .CO(n627), .S(n626) );
  ad01d0 U743 ( .A(n644), .B(n627), .CI(n646), .CO(n649), .S(n648) );
  xn02d1 U744 ( .A1(n930), .A2(n862), .ZN(product[7]) );
  aor21d1 U745 ( .B1(n774), .B2(n931), .A(n777), .Z(n930) );
  ad01d0 U746 ( .A(n514), .B(n491), .CI(n516), .CO(n523), .S(n522) );
  ad01d0 U747 ( .A(n488), .B(n490), .CI(n492), .CO(n497), .S(n496) );
  ad01d0 U748 ( .A(n521), .B(n546), .CI(n523), .CO(n553), .S(n552) );
  ad01d0 U749 ( .A(n443), .B(n464), .CI(n445), .CO(n471), .S(n470) );
  ad01d0 U750 ( .A(n493), .B(n518), .CI(n495), .CO(n525), .S(n524) );
  ad01d0 U751 ( .A(n404), .B(n389), .CI(n406), .CO(n409), .S(n408) );
  ad01d0 U752 ( .A(n424), .B(n407), .CI(n426), .CO(n429), .S(n428) );
  ad01d0 U753 ( .A(n359), .B(n370), .CI(n372), .CO(n375), .S(n374) );
  ad01d0 U754 ( .A(n347), .B(n356), .CI(n358), .CO(n361), .S(n360) );
  ad01d0 U755 ( .A(n373), .B(n386), .CI(n388), .CO(n391), .S(n390) );
  ad01d0 U756 ( .A(n400), .B(n387), .CI(n402), .CO(n407), .S(n406) );
  ad01d0 U757 ( .A(n442), .B(n444), .CI(n425), .CO(n449), .S(n448) );
  ad01d0 U758 ( .A(n420), .B(n405), .CI(n422), .CO(n427), .S(n426) );
  ad01d0 U759 ( .A(n519), .B(n542), .CI(n544), .CO(n551), .S(n550) );
  ad01d0 U760 ( .A(n466), .B(n447), .CI(n468), .CO(n473), .S(n472) );
  ad01d0 U761 ( .A(n469), .B(n471), .CI(n494), .CO(n499), .S(n498) );
  ad01d0 U762 ( .A(n548), .B(n525), .CI(n550), .CO(n555), .S(n554) );
  ad01d0 U763 ( .A(n520), .B(n522), .CI(n497), .CO(n527), .S(n526) );
  or02d1 U764 ( .A1(n348), .A2(n339), .Z(n931) );
  or02d1 U765 ( .A1(n360), .A2(n349), .Z(n932) );
  or02d1 U766 ( .A1(n338), .A2(n331), .Z(n933) );
  aoi21d1 U767 ( .B1(n934), .B2(n760), .A(n763), .ZN(n765) );
  inv0d1 U768 ( .I(n761), .ZN(n763) );
  ad01d0 U769 ( .A(n547), .B(n568), .CI(n570), .CO(n577), .S(n576) );
  ad01d0 U770 ( .A(n571), .B(n573), .CI(n594), .CO(n601), .S(n600) );
  ad01d0 U771 ( .A(n595), .B(n597), .CI(n616), .CO(n623), .S(n622) );
  ad01d0 U772 ( .A(n572), .B(n549), .CI(n574), .CO(n579), .S(n578) );
  ad01d0 U773 ( .A(n596), .B(n575), .CI(n598), .CO(n603), .S(n602) );
  ad01d0 U774 ( .A(n618), .B(n620), .CI(n599), .CO(n625), .S(n624) );
  ad01d0 U775 ( .A(n662), .B(n647), .CI(n664), .CO(n667), .S(n666) );
  ad01d0 U776 ( .A(n678), .B(n665), .CI(n680), .CO(n683), .S(n682) );
  ad01d0 U777 ( .A(n692), .B(n681), .CI(n694), .CO(n697), .S(n696) );
  ad01d0 U778 ( .A(n638), .B(n621), .CI(n640), .CO(n645), .S(n644) );
  ad01d0 U779 ( .A(n623), .B(n642), .CI(n625), .CO(n647), .S(n646) );
  ad01d0 U780 ( .A(n660), .B(n643), .CI(n645), .CO(n665), .S(n664) );
  ad01d0 U781 ( .A(n661), .B(n676), .CI(n663), .CO(n681), .S(n680) );
  ad01d0 U782 ( .A(n677), .B(n690), .CI(n679), .CO(n695), .S(n694) );
  ad01d0 U783 ( .A(n704), .B(n695), .CI(n706), .CO(n709), .S(n708) );
  ad01d0 U784 ( .A(n714), .B(n707), .CI(n716), .CO(n719), .S(n718) );
  ad01d0 U785 ( .A(n715), .B(n724), .CI(n717), .CO(n727), .S(n726) );
  inv0d1 U786 ( .I(n767), .ZN(n743) );
  inv0d1 U787 ( .I(n759), .ZN(n741) );
  ad01d0 U788 ( .A(n435), .B(n437), .CI(n460), .CO(n465), .S(n464) );
  ad01d0 U789 ( .A(n432), .B(n419), .CI(n438), .CO(n445), .S(n444) );
  ad01d0 U790 ( .A(n506), .B(n508), .CI(n504), .CO(n519), .S(n518) );
  ad01d0 U791 ( .A(n509), .B(n505), .CI(n511), .CO(n543), .S(n542) );
  ad01d0 U792 ( .A(n455), .B(n484), .CI(n482), .CO(n491), .S(n490) );
  ad01d0 U793 ( .A(n341), .B(n350), .CI(n343), .CO(n357), .S(n356) );
  ad01d0 U794 ( .A(n534), .B(n532), .CI(n513), .CO(n547), .S(n546) );
  ad01d0 U795 ( .A(n415), .B(n436), .CI(n434), .CO(n443), .S(n442) );
  ad01d0 U796 ( .A(n502), .B(n483), .CI(n479), .CO(n515), .S(n514) );
  ad01d0 U797 ( .A(n459), .B(n461), .CI(n457), .CO(n489), .S(n488) );
  ad01d0 U798 ( .A(n515), .B(n540), .CI(n517), .CO(n549), .S(n548) );
  ad01d0 U799 ( .A(n487), .B(n512), .CI(n489), .CO(n521), .S(n520) );
  ad01d0 U800 ( .A(n353), .B(n355), .CI(n366), .CO(n371), .S(n370) );
  ad01d0 U801 ( .A(n380), .B(n378), .CI(n369), .CO(n387), .S(n386) );
  ad01d0 U802 ( .A(n394), .B(n383), .CI(n385), .CO(n405), .S(n404) );
  ad01d0 U803 ( .A(n377), .B(n392), .CI(n379), .CO(n401), .S(n400) );
  ad01d0 U804 ( .A(n337), .B(n344), .CI(n346), .CO(n349), .S(n348) );
  ad01d0 U805 ( .A(n329), .B(n334), .CI(n336), .CO(n339), .S(n338) );
  ad01d0 U806 ( .A(n323), .B(n326), .CI(n328), .CO(n331), .S(n330) );
  ad01d0 U807 ( .A(n340), .B(n335), .CI(n342), .CO(n347), .S(n346) );
  ad01d0 U808 ( .A(n376), .B(n365), .CI(n367), .CO(n385), .S(n384) );
  ad01d0 U809 ( .A(n431), .B(n452), .CI(n433), .CO(n463), .S(n462) );
  ad01d0 U810 ( .A(n382), .B(n371), .CI(n384), .CO(n389), .S(n388) );
  ad01d0 U811 ( .A(n486), .B(n465), .CI(n467), .CO(n495), .S(n494) );
  ad01d0 U812 ( .A(n507), .B(n538), .CI(n536), .CO(n545), .S(n544) );
  ad01d0 U813 ( .A(n478), .B(n480), .CI(n463), .CO(n493), .S(n492) );
  ad01d0 U814 ( .A(n481), .B(n485), .CI(n510), .CO(n517), .S(n516) );
  ad01d0 U815 ( .A(n456), .B(n441), .CI(n462), .CO(n469), .S(n468) );
  ad01d0 U816 ( .A(n364), .B(n357), .CI(n368), .CO(n373), .S(n372) );
  ad01d0 U817 ( .A(n354), .B(n352), .CI(n345), .CO(n359), .S(n358) );
  ad01d0 U818 ( .A(n381), .B(n398), .CI(n396), .CO(n403), .S(n402) );
  ad01d0 U819 ( .A(n458), .B(n454), .CI(n439), .CO(n467), .S(n466) );
  ad01d0 U820 ( .A(n401), .B(n418), .CI(n403), .CO(n425), .S(n424) );
  ad01d0 U821 ( .A(n738), .B(n737), .CI(n853), .CO(n854), .S(product[29]) );
  or02d1 U822 ( .A1(n324), .A2(n322), .Z(n934) );
  ad01d0 U823 ( .A(n537), .B(n533), .CI(n539), .CO(n569), .S(n568) );
  ad01d0 U824 ( .A(n610), .B(n608), .CI(n593), .CO(n621), .S(n620) );
  ad01d0 U825 ( .A(n558), .B(n560), .CI(n541), .CO(n573), .S(n572) );
  ad01d0 U826 ( .A(n588), .B(n584), .CI(n567), .CO(n597), .S(n596) );
  ad01d0 U827 ( .A(n566), .B(n543), .CI(n545), .CO(n575), .S(n574) );
  ad01d0 U828 ( .A(n535), .B(n564), .CI(n562), .CO(n571), .S(n570) );
  ad01d0 U829 ( .A(n586), .B(n569), .CI(n592), .CO(n599), .S(n598) );
  ad01d0 U830 ( .A(n563), .B(n565), .CI(n590), .CO(n595), .S(n594) );
  ad01d0 U831 ( .A(n585), .B(n591), .CI(n589), .CO(n617), .S(n616) );
  ad01d0 U832 ( .A(n617), .B(n636), .CI(n619), .CO(n643), .S(n642) );
  ad01d0 U833 ( .A(n672), .B(n668), .CI(n670), .CO(n677), .S(n676) );
  ad01d0 U834 ( .A(n587), .B(n614), .CI(n612), .CO(n619), .S(n618) );
  ad01d0 U835 ( .A(n611), .B(n615), .CI(n613), .CO(n639), .S(n638) );
  ad01d0 U836 ( .A(n656), .B(n641), .CI(n658), .CO(n663), .S(n662) );
  ad01d0 U837 ( .A(n650), .B(n637), .CI(n639), .CO(n661), .S(n660) );
  ad01d0 U838 ( .A(n657), .B(n659), .CI(n674), .CO(n679), .S(n678) );
  ad01d0 U839 ( .A(n634), .B(n630), .CI(n632), .CO(n641), .S(n640) );
  ad01d0 U840 ( .A(n635), .B(n654), .CI(n652), .CO(n659), .S(n658) );
  ad01d0 U841 ( .A(n651), .B(n655), .CI(n653), .CO(n675), .S(n674) );
  ad01d0 U842 ( .A(n671), .B(n673), .CI(n686), .CO(n691), .S(n690) );
  ad01d0 U843 ( .A(n684), .B(n675), .CI(n688), .CO(n693), .S(n692) );
  ad01d0 U844 ( .A(n700), .B(n698), .CI(n689), .CO(n705), .S(n704) );
  ad01d0 U845 ( .A(n691), .B(n702), .CI(n693), .CO(n707), .S(n706) );
  ad01d0 U846 ( .A(n710), .B(n703), .CI(n705), .CO(n717), .S(n716) );
  ad01d0 U847 ( .A(n713), .B(n720), .CI(n722), .CO(n725), .S(n724) );
  ad01d0 U848 ( .A(n699), .B(n701), .CI(n712), .CO(n715), .S(n714) );
  ad01d0 U849 ( .A(n723), .B(n730), .CI(n725), .CO(n733), .S(n732) );
  ad01d0 U850 ( .A(n729), .B(n734), .CI(n731), .CO(n737), .S(n736) );
  an02d1 U851 ( .A1(n909), .A2(n756), .Z(product[1]) );
  ad01d0 U852 ( .A(n70), .B(n130), .CI(n85), .CO(n343), .S(n342) );
  ad01d0 U853 ( .A(n69), .B(n114), .CI(n99), .CO(n335), .S(n334) );
  ad01d0 U854 ( .A(n104), .B(n149), .CI(n119), .CO(n399), .S(n398) );
  ad01d0 U855 ( .A(n73), .B(n178), .CI(n88), .CO(n379), .S(n378) );
  ad01d0 U856 ( .A(n71), .B(n146), .CI(n86), .CO(n353), .S(n352) );
  ad01d0 U857 ( .A(n72), .B(n162), .CI(n87), .CO(n365), .S(n364) );
  ad01d0 U858 ( .A(n122), .B(n152), .CI(n137), .CO(n461), .S(n460) );
  ad01d0 U859 ( .A(n121), .B(n196), .CI(n181), .CO(n437), .S(n436) );
  ad01d0 U860 ( .A(n77), .B(n242), .CI(n92), .CO(n455), .S(n454) );
  ad01d0 U861 ( .A(n76), .B(n226), .CI(n211), .CO(n433), .S(n432) );
  ad01d0 U862 ( .A(n165), .B(n195), .CI(n180), .CO(n415), .S(n414) );
  ad01d0 U863 ( .A(n75), .B(n210), .CI(n90), .CO(n413), .S(n412) );
  ad01d0 U864 ( .A(n155), .B(n230), .CI(n185), .CO(n539), .S(n538) );
  ad01d0 U865 ( .A(n275), .B(n260), .CI(n245), .CO(n537), .S(n536) );
  ad01d0 U866 ( .A(n229), .B(n259), .CI(n244), .CO(n509), .S(n508) );
  ad01d0 U867 ( .A(n79), .B(n274), .CI(n94), .CO(n505), .S(n504) );
  ad01d0 U868 ( .A(n139), .B(n214), .CI(n184), .CO(n511), .S(n510) );
  ad01d0 U869 ( .A(n168), .B(n228), .CI(n93), .CO(n481), .S(n480) );
  ad01d0 U870 ( .A(n123), .B(n198), .CI(n153), .CO(n485), .S(n484) );
  ad01d0 U871 ( .A(n183), .B(n108), .CI(n213), .CO(n483), .S(n482) );
  ad01d0 U872 ( .A(n200), .B(n95), .CI(n110), .CO(n533), .S(n532) );
  ad01d0 U873 ( .A(n169), .B(n154), .CI(n477), .CO(n513), .S(n512) );
  ad01d0 U874 ( .A(n170), .B(n503), .CI(n530), .CO(n541), .S(n540) );
  ad01d0 U875 ( .A(n101), .B(n131), .CI(n116), .CO(n355), .S(n354) );
  ad01d0 U876 ( .A(n107), .B(n197), .CI(n167), .CO(n459), .S(n458) );
  ad01d0 U877 ( .A(n103), .B(n118), .CI(n363), .CO(n383), .S(n382) );
  ad01d0 U878 ( .A(n105), .B(n150), .CI(n135), .CO(n417), .S(n416) );
  ad01d0 U879 ( .A(n199), .B(n109), .CI(n124), .CO(n507), .S(n506) );
  ad01d0 U880 ( .A(n78), .B(n258), .CI(n243), .CO(n479), .S(n478) );
  ad01d0 U881 ( .A(n182), .B(n227), .CI(n212), .CO(n457), .S(n456) );
  ad01d0 U882 ( .A(n215), .B(n125), .CI(n140), .CO(n535), .S(n534) );
  ad01d0 U883 ( .A(n138), .B(n453), .CI(n476), .CO(n487), .S(n486) );
  ad01d0 U884 ( .A(n120), .B(n393), .CI(n410), .CO(n419), .S(n418) );
  ad01d0 U885 ( .A(n148), .B(n163), .CI(n133), .CO(n381), .S(n380) );
  ad01d0 U886 ( .A(n166), .B(n91), .CI(n106), .CO(n435), .S(n434) );
  ad01d0 U887 ( .A(n74), .B(n194), .CI(n179), .CO(n395), .S(n394) );
  ad01d0 U888 ( .A(n67), .B(n82), .CI(n321), .CO(n325), .S(n324) );
  ad01d0 U889 ( .A(n84), .B(n327), .CI(n332), .CO(n337), .S(n336) );
  ad01d0 U890 ( .A(n68), .B(n98), .CI(n83), .CO(n329), .S(n328) );
  ad01d0 U891 ( .A(n134), .B(n89), .CI(n164), .CO(n397), .S(n396) );
  ad01d0 U892 ( .A(n117), .B(n351), .CI(n362), .CO(n369), .S(n368) );
  ad01d0 U893 ( .A(n132), .B(n102), .CI(n147), .CO(n367), .S(n366) );
  ad01d0 U894 ( .A(n136), .B(n151), .CI(n411), .CO(n439), .S(n438) );
  ad01d0 U895 ( .A(n100), .B(n115), .CI(n333), .CO(n345), .S(n344) );
  ad01d0 U896 ( .A(n319), .B(n739), .CI(n854), .CO(product[31]), .S(
        product[30]) );
  ad01d0 U897 ( .A(n201), .B(n126), .CI(n276), .CO(n561), .S(n560) );
  ad01d0 U898 ( .A(n141), .B(n261), .CI(n156), .CO(n563), .S(n562) );
  ad01d0 U899 ( .A(n171), .B(n246), .CI(n231), .CO(n565), .S(n564) );
  ad01d0 U900 ( .A(n127), .B(n307), .CI(n142), .CO(n585), .S(n584) );
  ad01d0 U901 ( .A(n187), .B(n232), .CI(n217), .CO(n591), .S(n590) );
  ad01d0 U902 ( .A(n111), .B(n306), .CI(n291), .CO(n559), .S(n558) );
  ad01d0 U903 ( .A(n186), .B(n216), .CI(n531), .CO(n567), .S(n566) );
  ad01d0 U904 ( .A(n157), .B(n292), .CI(n277), .CO(n587), .S(n586) );
  ad01d0 U905 ( .A(n247), .B(n172), .CI(n262), .CO(n589), .S(n588) );
  ad01d0 U906 ( .A(n202), .B(n559), .CI(n561), .CO(n593), .S(n592) );
  ad01d0 U907 ( .A(n143), .B(n308), .CI(n293), .CO(n609), .S(n608) );
  ad01d0 U908 ( .A(n188), .B(n218), .CI(n203), .CO(n615), .S(n614) );
  ad01d0 U909 ( .A(n159), .B(n309), .CI(n294), .CO(n631), .S(n630) );
  ad01d0 U910 ( .A(n174), .B(n279), .CI(n264), .CO(n633), .S(n632) );
  ad01d0 U911 ( .A(n220), .B(n265), .CI(n250), .CO(n655), .S(n654) );
  ad01d0 U912 ( .A(n190), .B(n280), .CI(n205), .CO(n653), .S(n652) );
  ad01d0 U913 ( .A(n191), .B(n311), .CI(n296), .CO(n669), .S(n668) );
  ad01d0 U914 ( .A(n189), .B(n204), .CI(n609), .CO(n637), .S(n636) );
  ad01d0 U915 ( .A(n158), .B(n278), .CI(n263), .CO(n611), .S(n610) );
  ad01d0 U916 ( .A(n219), .B(n249), .CI(n234), .CO(n635), .S(n634) );
  ad01d0 U917 ( .A(n175), .B(n310), .CI(n295), .CO(n651), .S(n650) );
  ad01d0 U918 ( .A(n236), .B(n266), .CI(n251), .CO(n673), .S(n672) );
  ad01d0 U919 ( .A(n235), .B(n631), .CI(n633), .CO(n657), .S(n656) );
  ad01d0 U920 ( .A(n248), .B(n173), .CI(n233), .CO(n613), .S(n612) );
  ad01d0 U921 ( .A(n206), .B(n281), .CI(n221), .CO(n671), .S(n670) );
  ad01d0 U922 ( .A(n223), .B(n313), .CI(n298), .CO(n699), .S(n698) );
  ad01d0 U923 ( .A(n268), .B(n685), .CI(n687), .CO(n703), .S(n702) );
  ad01d0 U924 ( .A(n283), .B(n238), .CI(n253), .CO(n701), .S(n700) );
  ad01d0 U925 ( .A(n207), .B(n312), .CI(n297), .CO(n685), .S(n684) );
  ad01d0 U926 ( .A(n237), .B(n252), .CI(n669), .CO(n689), .S(n688) );
  ad01d0 U927 ( .A(n222), .B(n282), .CI(n267), .CO(n687), .S(n686) );
  ad01d0 U928 ( .A(n255), .B(n315), .CI(n300), .CO(n721), .S(n720) );
  ad01d0 U929 ( .A(n286), .B(n721), .CI(n728), .CO(n731), .S(n730) );
  ad01d0 U930 ( .A(n239), .B(n314), .CI(n299), .CO(n711), .S(n710) );
  ad01d0 U931 ( .A(n270), .B(n285), .CI(n711), .CO(n723), .S(n722) );
  ad01d0 U932 ( .A(n284), .B(n269), .CI(n254), .CO(n713), .S(n712) );
  ad01d0 U933 ( .A(n271), .B(n316), .CI(n301), .CO(n729), .S(n728) );
  ad01d0 U934 ( .A(n287), .B(n317), .CI(n302), .CO(n735), .S(n734) );
  ad01d0 U935 ( .A(n303), .B(n318), .CI(n735), .CO(n739), .S(n738) );
  inv0d1 U936 ( .I(a[0]), .ZN(n32) );
  inv0d1 U937 ( .I(a[3]), .ZN(n35) );
  inv0d1 U938 ( .I(a[4]), .ZN(n36) );
  inv0d1 U939 ( .I(a[6]), .ZN(n38) );
  inv0d1 U940 ( .I(a[7]), .ZN(n39) );
  inv0d1 U941 ( .I(a[8]), .ZN(n40) );
  inv0d1 U942 ( .I(a[10]), .ZN(n42) );
  inv0d1 U943 ( .I(a[13]), .ZN(n45) );
  inv0d1 U944 ( .I(a[14]), .ZN(n46) );
  inv0d1 U945 ( .I(a[15]), .ZN(n47) );
  inv0d1 U946 ( .I(b[0]), .ZN(n48) );
  inv0d1 U947 ( .I(b[1]), .ZN(n49) );
  inv0d1 U948 ( .I(b[3]), .ZN(n51) );
  inv0d1 U949 ( .I(b[4]), .ZN(n52) );
  inv0d1 U950 ( .I(b[5]), .ZN(n53) );
  inv0d1 U951 ( .I(b[7]), .ZN(n55) );
  inv0d1 U952 ( .I(b[8]), .ZN(n56) );
  inv0d1 U953 ( .I(b[10]), .ZN(n58) );
  inv0d1 U954 ( .I(b[12]), .ZN(n60) );
  inv0d1 U955 ( .I(b[13]), .ZN(n61) );
  inv0d1 U956 ( .I(b[14]), .ZN(n62) );
  inv0d1 U957 ( .I(b[15]), .ZN(n63) );
endmodule


module BLENDER_DW_mult_uns_6 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n741, n743, n747, n748, n753, n756, n758, n759, n760, n761, n763,
         n765, n766, n767, n768, n769, n771, n773, n774, n775, n777, n780,
         n782, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n799, n802, n804, n806, n807, n808, n809,
         n812, n813, n814, n815, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n832, n835, n837, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937;

  nr02d0 U33 ( .A1(n48), .A2(n925), .ZN(product[0]) );
  nr02d0 U34 ( .A1(n49), .A2(n32), .ZN(n65) );
  nr02d0 U35 ( .A1(n50), .A2(n925), .ZN(n66) );
  nr02d0 U36 ( .A1(n51), .A2(n925), .ZN(n67) );
  nr02d0 U37 ( .A1(n52), .A2(n32), .ZN(n68) );
  nr02d0 U38 ( .A1(n53), .A2(n32), .ZN(n69) );
  nr02d0 U39 ( .A1(n54), .A2(n32), .ZN(n70) );
  nr02d0 U40 ( .A1(n55), .A2(n32), .ZN(n71) );
  nr02d0 U41 ( .A1(n56), .A2(n925), .ZN(n72) );
  nr02d0 U42 ( .A1(n57), .A2(n925), .ZN(n73) );
  nr02d0 U43 ( .A1(n58), .A2(n32), .ZN(n74) );
  nr02d0 U44 ( .A1(n59), .A2(n32), .ZN(n75) );
  nr02d0 U45 ( .A1(n60), .A2(n925), .ZN(n76) );
  nr02d0 U46 ( .A1(n61), .A2(n925), .ZN(n77) );
  nr02d0 U47 ( .A1(n62), .A2(n925), .ZN(n78) );
  nr02d0 U48 ( .A1(n63), .A2(n32), .ZN(n79) );
  nr02d0 U49 ( .A1(n48), .A2(n33), .ZN(n80) );
  nr02d0 U50 ( .A1(n49), .A2(n33), .ZN(n81) );
  nr02d0 U51 ( .A1(n50), .A2(n33), .ZN(n82) );
  nr02d0 U52 ( .A1(n51), .A2(n33), .ZN(n83) );
  nr02d0 U53 ( .A1(n52), .A2(n33), .ZN(n84) );
  nr02d0 U54 ( .A1(n53), .A2(n33), .ZN(n85) );
  nr02d0 U55 ( .A1(n54), .A2(n33), .ZN(n86) );
  nr02d0 U56 ( .A1(n55), .A2(n33), .ZN(n87) );
  nr02d0 U57 ( .A1(n56), .A2(n33), .ZN(n88) );
  nr02d0 U58 ( .A1(n57), .A2(n33), .ZN(n89) );
  nr02d0 U59 ( .A1(n58), .A2(n33), .ZN(n90) );
  nr02d0 U60 ( .A1(n59), .A2(n33), .ZN(n91) );
  nr02d0 U61 ( .A1(n60), .A2(n33), .ZN(n92) );
  nr02d0 U62 ( .A1(n61), .A2(n33), .ZN(n93) );
  nr02d0 U63 ( .A1(n62), .A2(n33), .ZN(n94) );
  nr02d0 U64 ( .A1(n63), .A2(n33), .ZN(n95) );
  nr02d0 U65 ( .A1(n48), .A2(n34), .ZN(n96) );
  nr02d0 U66 ( .A1(n49), .A2(n34), .ZN(n97) );
  nr02d0 U67 ( .A1(n50), .A2(n34), .ZN(n98) );
  nr02d0 U68 ( .A1(n51), .A2(n34), .ZN(n99) );
  nr02d0 U69 ( .A1(n52), .A2(n34), .ZN(n100) );
  nr02d0 U71 ( .A1(n54), .A2(n34), .ZN(n102) );
  nr02d0 U72 ( .A1(n55), .A2(n34), .ZN(n103) );
  nr02d0 U73 ( .A1(n56), .A2(n34), .ZN(n104) );
  nr02d0 U74 ( .A1(n57), .A2(n34), .ZN(n105) );
  nr02d0 U75 ( .A1(n58), .A2(n34), .ZN(n106) );
  nr02d0 U76 ( .A1(n59), .A2(n34), .ZN(n107) );
  nr02d0 U77 ( .A1(n60), .A2(n34), .ZN(n108) );
  nr02d0 U78 ( .A1(n61), .A2(n34), .ZN(n109) );
  nr02d0 U79 ( .A1(n62), .A2(n34), .ZN(n110) );
  nr02d0 U80 ( .A1(n63), .A2(n34), .ZN(n111) );
  nr02d0 U81 ( .A1(n48), .A2(n35), .ZN(n112) );
  nr02d0 U82 ( .A1(n49), .A2(n35), .ZN(n113) );
  nr02d0 U83 ( .A1(n50), .A2(n35), .ZN(n114) );
  nr02d0 U84 ( .A1(n51), .A2(n35), .ZN(n115) );
  nr02d0 U85 ( .A1(n52), .A2(n35), .ZN(n116) );
  nr02d0 U86 ( .A1(n53), .A2(n35), .ZN(n117) );
  nr02d0 U87 ( .A1(n54), .A2(n35), .ZN(n118) );
  nr02d0 U88 ( .A1(n55), .A2(n35), .ZN(n119) );
  nr02d0 U89 ( .A1(n56), .A2(n35), .ZN(n120) );
  nr02d0 U90 ( .A1(n57), .A2(n35), .ZN(n121) );
  nr02d0 U91 ( .A1(n58), .A2(n35), .ZN(n122) );
  nr02d0 U92 ( .A1(n59), .A2(n35), .ZN(n123) );
  nr02d0 U93 ( .A1(n60), .A2(n35), .ZN(n124) );
  nr02d0 U94 ( .A1(n61), .A2(n35), .ZN(n125) );
  nr02d0 U95 ( .A1(n62), .A2(n35), .ZN(n126) );
  nr02d0 U96 ( .A1(n63), .A2(n35), .ZN(n127) );
  nr02d0 U97 ( .A1(n48), .A2(n36), .ZN(n128) );
  nr02d0 U98 ( .A1(n49), .A2(n36), .ZN(n129) );
  nr02d0 U99 ( .A1(n50), .A2(n36), .ZN(n130) );
  nr02d0 U100 ( .A1(n51), .A2(n36), .ZN(n131) );
  nr02d0 U101 ( .A1(n52), .A2(n36), .ZN(n132) );
  nr02d0 U102 ( .A1(n53), .A2(n36), .ZN(n133) );
  nr02d0 U104 ( .A1(n55), .A2(n36), .ZN(n135) );
  nr02d0 U105 ( .A1(n56), .A2(n36), .ZN(n136) );
  nr02d0 U106 ( .A1(n57), .A2(n36), .ZN(n137) );
  nr02d0 U107 ( .A1(n58), .A2(n36), .ZN(n138) );
  nr02d0 U108 ( .A1(n59), .A2(n36), .ZN(n139) );
  nr02d0 U109 ( .A1(n60), .A2(n36), .ZN(n140) );
  nr02d0 U110 ( .A1(n61), .A2(n36), .ZN(n141) );
  nr02d0 U111 ( .A1(n62), .A2(n36), .ZN(n142) );
  nr02d0 U112 ( .A1(n63), .A2(n36), .ZN(n143) );
  nr02d0 U113 ( .A1(n48), .A2(n37), .ZN(n144) );
  nr02d0 U114 ( .A1(n49), .A2(n37), .ZN(n145) );
  nr02d0 U115 ( .A1(n50), .A2(n37), .ZN(n146) );
  nr02d0 U117 ( .A1(n52), .A2(n37), .ZN(n148) );
  nr02d0 U118 ( .A1(n53), .A2(n37), .ZN(n149) );
  nr02d0 U119 ( .A1(n54), .A2(n37), .ZN(n150) );
  nr02d0 U120 ( .A1(n55), .A2(n37), .ZN(n151) );
  nr02d0 U121 ( .A1(n56), .A2(n37), .ZN(n152) );
  nr02d0 U122 ( .A1(n57), .A2(n37), .ZN(n153) );
  nr02d0 U123 ( .A1(n58), .A2(n37), .ZN(n154) );
  nr02d0 U124 ( .A1(n59), .A2(n37), .ZN(n155) );
  nr02d0 U125 ( .A1(n60), .A2(n37), .ZN(n156) );
  nr02d0 U126 ( .A1(n61), .A2(n37), .ZN(n157) );
  nr02d0 U127 ( .A1(n62), .A2(n37), .ZN(n158) );
  nr02d0 U128 ( .A1(n63), .A2(n37), .ZN(n159) );
  nr02d0 U129 ( .A1(n48), .A2(n38), .ZN(n160) );
  nr02d0 U130 ( .A1(n49), .A2(n38), .ZN(n161) );
  nr02d0 U131 ( .A1(n50), .A2(n38), .ZN(n162) );
  nr02d0 U132 ( .A1(n51), .A2(n38), .ZN(n163) );
  nr02d0 U133 ( .A1(n52), .A2(n38), .ZN(n164) );
  nr02d0 U134 ( .A1(n53), .A2(n38), .ZN(n165) );
  nr02d0 U136 ( .A1(n55), .A2(n38), .ZN(n167) );
  nr02d0 U137 ( .A1(n56), .A2(n916), .ZN(n168) );
  nr02d0 U138 ( .A1(n57), .A2(n916), .ZN(n169) );
  nr02d0 U139 ( .A1(n58), .A2(n916), .ZN(n170) );
  nr02d0 U140 ( .A1(n59), .A2(n916), .ZN(n171) );
  nr02d0 U141 ( .A1(n60), .A2(n916), .ZN(n172) );
  nr02d0 U142 ( .A1(n61), .A2(n916), .ZN(n173) );
  nr02d0 U143 ( .A1(n62), .A2(n916), .ZN(n174) );
  nr02d0 U144 ( .A1(n63), .A2(n916), .ZN(n175) );
  nr02d0 U145 ( .A1(n48), .A2(n39), .ZN(n176) );
  nr02d0 U146 ( .A1(n49), .A2(n39), .ZN(n177) );
  nr02d0 U147 ( .A1(n50), .A2(n39), .ZN(n178) );
  nr02d0 U148 ( .A1(n51), .A2(n39), .ZN(n179) );
  nr02d0 U149 ( .A1(n52), .A2(n39), .ZN(n180) );
  nr02d0 U150 ( .A1(n53), .A2(n39), .ZN(n181) );
  nr02d0 U151 ( .A1(n54), .A2(n39), .ZN(n182) );
  nr02d0 U152 ( .A1(n55), .A2(n39), .ZN(n183) );
  nr02d0 U153 ( .A1(n56), .A2(n39), .ZN(n184) );
  nr02d0 U154 ( .A1(n57), .A2(n39), .ZN(n185) );
  nr02d0 U155 ( .A1(n58), .A2(n39), .ZN(n186) );
  nr02d0 U156 ( .A1(n59), .A2(n39), .ZN(n187) );
  nr02d0 U157 ( .A1(n60), .A2(n39), .ZN(n188) );
  nr02d0 U158 ( .A1(n61), .A2(n39), .ZN(n189) );
  nr02d0 U159 ( .A1(n62), .A2(n39), .ZN(n190) );
  nr02d0 U160 ( .A1(n63), .A2(n39), .ZN(n191) );
  nr02d0 U161 ( .A1(n48), .A2(n40), .ZN(n192) );
  nr02d0 U162 ( .A1(n49), .A2(n40), .ZN(n193) );
  nr02d0 U163 ( .A1(n50), .A2(n40), .ZN(n194) );
  nr02d0 U164 ( .A1(n51), .A2(n40), .ZN(n195) );
  nr02d0 U165 ( .A1(n52), .A2(n40), .ZN(n196) );
  nr02d0 U166 ( .A1(n53), .A2(n40), .ZN(n197) );
  nr02d0 U167 ( .A1(n54), .A2(n40), .ZN(n198) );
  nr02d0 U168 ( .A1(n55), .A2(n40), .ZN(n199) );
  nr02d0 U169 ( .A1(n56), .A2(n915), .ZN(n200) );
  nr02d0 U170 ( .A1(n57), .A2(n915), .ZN(n201) );
  nr02d0 U171 ( .A1(n58), .A2(n915), .ZN(n202) );
  nr02d0 U172 ( .A1(n59), .A2(n915), .ZN(n203) );
  nr02d0 U173 ( .A1(n911), .A2(n915), .ZN(n204) );
  nr02d0 U174 ( .A1(n61), .A2(n915), .ZN(n205) );
  nr02d0 U175 ( .A1(n62), .A2(n915), .ZN(n206) );
  nr02d0 U176 ( .A1(n63), .A2(n915), .ZN(n207) );
  nr02d0 U177 ( .A1(n48), .A2(n41), .ZN(n208) );
  nr02d0 U178 ( .A1(n49), .A2(n41), .ZN(n209) );
  nr02d0 U179 ( .A1(n50), .A2(n41), .ZN(n210) );
  nr02d0 U180 ( .A1(n51), .A2(n41), .ZN(n211) );
  nr02d0 U181 ( .A1(n52), .A2(n41), .ZN(n212) );
  nr02d0 U182 ( .A1(n53), .A2(n41), .ZN(n213) );
  nr02d0 U183 ( .A1(n54), .A2(n41), .ZN(n214) );
  nr02d0 U184 ( .A1(n55), .A2(n41), .ZN(n215) );
  nr02d0 U185 ( .A1(n56), .A2(n41), .ZN(n216) );
  nr02d0 U186 ( .A1(n57), .A2(n41), .ZN(n217) );
  nr02d0 U187 ( .A1(n58), .A2(n41), .ZN(n218) );
  nr02d0 U188 ( .A1(n59), .A2(n41), .ZN(n219) );
  nr02d0 U189 ( .A1(n911), .A2(n41), .ZN(n220) );
  nr02d0 U190 ( .A1(n61), .A2(n41), .ZN(n221) );
  nr02d0 U191 ( .A1(n62), .A2(n41), .ZN(n222) );
  nr02d0 U192 ( .A1(n63), .A2(n41), .ZN(n223) );
  nr02d0 U193 ( .A1(n48), .A2(n42), .ZN(n224) );
  nr02d0 U194 ( .A1(n49), .A2(n42), .ZN(n225) );
  nr02d0 U195 ( .A1(n50), .A2(n42), .ZN(n226) );
  nr02d0 U196 ( .A1(n51), .A2(n42), .ZN(n227) );
  nr02d0 U197 ( .A1(n52), .A2(n42), .ZN(n228) );
  nr02d0 U198 ( .A1(n53), .A2(n42), .ZN(n229) );
  nr02d0 U199 ( .A1(n54), .A2(n42), .ZN(n230) );
  nr02d0 U200 ( .A1(n55), .A2(n42), .ZN(n231) );
  nr02d0 U201 ( .A1(n56), .A2(n913), .ZN(n232) );
  nr02d0 U202 ( .A1(n57), .A2(n913), .ZN(n233) );
  nr02d0 U203 ( .A1(n58), .A2(n913), .ZN(n234) );
  nr02d0 U204 ( .A1(n59), .A2(n913), .ZN(n235) );
  nr02d0 U205 ( .A1(n911), .A2(n913), .ZN(n236) );
  nr02d0 U206 ( .A1(n61), .A2(n913), .ZN(n237) );
  nr02d0 U207 ( .A1(n62), .A2(n913), .ZN(n238) );
  nr02d0 U208 ( .A1(n63), .A2(n913), .ZN(n239) );
  nr02d0 U209 ( .A1(n48), .A2(n43), .ZN(n240) );
  nr02d0 U210 ( .A1(n49), .A2(n43), .ZN(n241) );
  nr02d0 U211 ( .A1(n50), .A2(n43), .ZN(n242) );
  nr02d0 U212 ( .A1(n51), .A2(n43), .ZN(n243) );
  nr02d0 U213 ( .A1(n52), .A2(n43), .ZN(n244) );
  nr02d0 U214 ( .A1(n53), .A2(n43), .ZN(n245) );
  nr02d0 U215 ( .A1(n54), .A2(n43), .ZN(n246) );
  nr02d0 U216 ( .A1(n55), .A2(n43), .ZN(n247) );
  nr02d0 U217 ( .A1(n56), .A2(n43), .ZN(n248) );
  nr02d0 U218 ( .A1(n57), .A2(n43), .ZN(n249) );
  nr02d0 U219 ( .A1(n58), .A2(n43), .ZN(n250) );
  nr02d0 U220 ( .A1(n59), .A2(n43), .ZN(n251) );
  nr02d0 U221 ( .A1(n911), .A2(n43), .ZN(n252) );
  nr02d0 U222 ( .A1(n61), .A2(n43), .ZN(n253) );
  nr02d0 U223 ( .A1(n62), .A2(n43), .ZN(n254) );
  nr02d0 U224 ( .A1(n63), .A2(n43), .ZN(n255) );
  nr02d0 U225 ( .A1(n48), .A2(n44), .ZN(n256) );
  nr02d0 U226 ( .A1(n49), .A2(n44), .ZN(n257) );
  nr02d0 U227 ( .A1(n50), .A2(n44), .ZN(n258) );
  nr02d0 U228 ( .A1(n51), .A2(n44), .ZN(n259) );
  nr02d0 U229 ( .A1(n52), .A2(n44), .ZN(n260) );
  nr02d0 U230 ( .A1(n53), .A2(n44), .ZN(n261) );
  nr02d0 U231 ( .A1(n54), .A2(n44), .ZN(n262) );
  nr02d0 U232 ( .A1(n55), .A2(n44), .ZN(n263) );
  nr02d0 U233 ( .A1(n56), .A2(n44), .ZN(n264) );
  nr02d0 U234 ( .A1(n57), .A2(n44), .ZN(n265) );
  nr02d0 U235 ( .A1(n58), .A2(n44), .ZN(n266) );
  nr02d0 U236 ( .A1(n59), .A2(n44), .ZN(n267) );
  nr02d0 U237 ( .A1(n911), .A2(n44), .ZN(n268) );
  nr02d0 U238 ( .A1(n61), .A2(n44), .ZN(n269) );
  nr02d0 U239 ( .A1(n62), .A2(n44), .ZN(n270) );
  nr02d0 U240 ( .A1(n63), .A2(n44), .ZN(n271) );
  nr02d0 U242 ( .A1(n49), .A2(n45), .ZN(n273) );
  nr02d0 U243 ( .A1(n50), .A2(n45), .ZN(n274) );
  nr02d0 U244 ( .A1(n51), .A2(n45), .ZN(n275) );
  nr02d0 U245 ( .A1(n52), .A2(n45), .ZN(n276) );
  nr02d0 U246 ( .A1(n53), .A2(n45), .ZN(n277) );
  nr02d0 U247 ( .A1(n54), .A2(n45), .ZN(n278) );
  nr02d0 U248 ( .A1(n55), .A2(n45), .ZN(n279) );
  nr02d0 U249 ( .A1(n56), .A2(n45), .ZN(n280) );
  nr02d0 U250 ( .A1(n57), .A2(n45), .ZN(n281) );
  nr02d0 U251 ( .A1(n58), .A2(n45), .ZN(n282) );
  nr02d0 U252 ( .A1(n59), .A2(n45), .ZN(n283) );
  nr02d0 U253 ( .A1(n911), .A2(n45), .ZN(n284) );
  nr02d0 U254 ( .A1(n61), .A2(n45), .ZN(n285) );
  nr02d0 U255 ( .A1(n62), .A2(n45), .ZN(n286) );
  nr02d0 U256 ( .A1(n63), .A2(n45), .ZN(n287) );
  nr02d0 U257 ( .A1(n48), .A2(n46), .ZN(n288) );
  nr02d0 U258 ( .A1(n49), .A2(n46), .ZN(n289) );
  nr02d0 U259 ( .A1(n50), .A2(n46), .ZN(n290) );
  nr02d0 U260 ( .A1(n51), .A2(n46), .ZN(n291) );
  nr02d0 U261 ( .A1(n52), .A2(n46), .ZN(n292) );
  nr02d0 U262 ( .A1(n53), .A2(n46), .ZN(n293) );
  nr02d0 U263 ( .A1(n54), .A2(n46), .ZN(n294) );
  nr02d0 U264 ( .A1(n55), .A2(n46), .ZN(n295) );
  nr02d0 U265 ( .A1(n56), .A2(n46), .ZN(n296) );
  nr02d0 U266 ( .A1(n57), .A2(n46), .ZN(n297) );
  nr02d0 U267 ( .A1(n58), .A2(n46), .ZN(n298) );
  nr02d0 U268 ( .A1(n59), .A2(n46), .ZN(n299) );
  nr02d0 U269 ( .A1(n911), .A2(n46), .ZN(n300) );
  nr02d0 U270 ( .A1(n61), .A2(n46), .ZN(n301) );
  nr02d0 U271 ( .A1(n62), .A2(n46), .ZN(n302) );
  nr02d0 U272 ( .A1(n63), .A2(n46), .ZN(n303) );
  nr02d0 U273 ( .A1(n48), .A2(n47), .ZN(n304) );
  nr02d0 U274 ( .A1(n49), .A2(n47), .ZN(n305) );
  nr02d0 U275 ( .A1(n50), .A2(n47), .ZN(n306) );
  nr02d0 U276 ( .A1(n51), .A2(n47), .ZN(n307) );
  nr02d0 U277 ( .A1(n52), .A2(n47), .ZN(n308) );
  nr02d0 U278 ( .A1(n53), .A2(n47), .ZN(n309) );
  nr02d0 U279 ( .A1(n54), .A2(n47), .ZN(n310) );
  nr02d0 U280 ( .A1(n55), .A2(n47), .ZN(n311) );
  nr02d0 U281 ( .A1(n56), .A2(n47), .ZN(n312) );
  nr02d0 U282 ( .A1(n57), .A2(n47), .ZN(n313) );
  nr02d0 U283 ( .A1(n58), .A2(n47), .ZN(n314) );
  nr02d0 U284 ( .A1(n59), .A2(n47), .ZN(n315) );
  nr02d0 U285 ( .A1(n911), .A2(n47), .ZN(n316) );
  nr02d0 U286 ( .A1(n61), .A2(n47), .ZN(n317) );
  nr02d0 U287 ( .A1(n62), .A2(n47), .ZN(n318) );
  nr02d0 U288 ( .A1(n63), .A2(n47), .ZN(n319) );
  ah01d0 U289 ( .A(n66), .B(n81), .CO(n321), .S(n320) );
  ah01d0 U290 ( .A(n97), .B(n112), .CO(n323), .S(n322) );
  ah01d0 U292 ( .A(n113), .B(n128), .CO(n327), .S(n326) );
  ah01d0 U295 ( .A(n129), .B(n144), .CO(n333), .S(n332) );
  ah01d0 U299 ( .A(n145), .B(n160), .CO(n341), .S(n340) );
  ah01d0 U304 ( .A(n161), .B(n176), .CO(n351), .S(n350) );
  ah01d0 U310 ( .A(n177), .B(n192), .CO(n363), .S(n362) );
  ah01d0 U317 ( .A(n193), .B(n208), .CO(n377), .S(n376) );
  ah01d0 U325 ( .A(n209), .B(n224), .CO(n393), .S(n392) );
  ah01d0 U334 ( .A(n225), .B(n240), .CO(n411), .S(n410) );
  ah01d0 U344 ( .A(n241), .B(n256), .CO(n431), .S(n430) );
  ah01d0 U367 ( .A(n273), .B(n288), .CO(n477), .S(n476) );
  ah01d0 U380 ( .A(n289), .B(n304), .CO(n503), .S(n502) );
  ah01d0 U394 ( .A(n290), .B(n305), .CO(n531), .S(n530) );
  nd02d1 U499 ( .A1(n65), .A2(n80), .ZN(n756) );
  nd02d1 U504 ( .A1(n320), .A2(n96), .ZN(n758) );
  nr02d0 U505 ( .A1(n320), .A2(n96), .ZN(n759) );
  nd02d1 U507 ( .A1(n741), .A2(n758), .ZN(n857) );
  oai21d1 U508 ( .B1(n759), .B2(n756), .A(n758), .ZN(n760) );
  xr02d1 U509 ( .A1(n857), .A2(n756), .Z(product[2]) );
  nd02d1 U510 ( .A1(n324), .A2(n322), .ZN(n761) );
  nd02d1 U513 ( .A1(n937), .A2(n761), .ZN(n858) );
  xn02d1 U517 ( .A1(n858), .A2(n760), .ZN(product[3]) );
  nd02d1 U518 ( .A1(n330), .A2(n325), .ZN(n766) );
  nr02d0 U519 ( .A1(n330), .A2(n325), .ZN(n767) );
  nd02d1 U521 ( .A1(n743), .A2(n766), .ZN(n859) );
  oai21d1 U522 ( .B1(n767), .B2(n765), .A(n766), .ZN(n768) );
  xr02d1 U523 ( .A1(n859), .A2(n765), .Z(product[4]) );
  nd02d1 U524 ( .A1(n338), .A2(n331), .ZN(n769) );
  nd02d1 U527 ( .A1(n936), .A2(n769), .ZN(n860) );
  xn02d1 U532 ( .A1(n860), .A2(n768), .ZN(product[5]) );
  nd02d1 U533 ( .A1(n348), .A2(n339), .ZN(n775) );
  nd02d1 U536 ( .A1(n934), .A2(n775), .ZN(n861) );
  xn02d1 U540 ( .A1(n861), .A2(n774), .ZN(product[6]) );
  nd02d1 U541 ( .A1(n360), .A2(n349), .ZN(n780) );
  nd02d1 U544 ( .A1(n935), .A2(n780), .ZN(n862) );
  nd02d1 U548 ( .A1(n935), .A2(n934), .ZN(n785) );
  oai21d1 U549 ( .B1(n785), .B2(n773), .A(n784), .ZN(n786) );
  nd02d1 U552 ( .A1(n374), .A2(n361), .ZN(n788) );
  nr02d0 U553 ( .A1(n374), .A2(n361), .ZN(n789) );
  nd02d1 U555 ( .A1(n747), .A2(n788), .ZN(n863) );
  oai21d1 U556 ( .B1(n787), .B2(n789), .A(n788), .ZN(n790) );
  xr02d1 U557 ( .A1(n787), .A2(n863), .Z(product[8]) );
  nd02d1 U558 ( .A1(n390), .A2(n375), .ZN(n791) );
  nr02d0 U559 ( .A1(n390), .A2(n375), .ZN(n792) );
  nd02d1 U561 ( .A1(n748), .A2(n791), .ZN(n864) );
  oai21d1 U562 ( .B1(n792), .B2(n788), .A(n791), .ZN(n793) );
  nr02d0 U563 ( .A1(n792), .A2(n789), .ZN(n794) );
  xn02d1 U566 ( .A1(n790), .A2(n864), .ZN(product[9]) );
  nd02d1 U567 ( .A1(n408), .A2(n391), .ZN(n797) );
  nd02d1 U570 ( .A1(n931), .A2(n797), .ZN(n865) );
  xn02d1 U574 ( .A1(n796), .A2(n865), .ZN(product[10]) );
  nd02d1 U575 ( .A1(n428), .A2(n409), .ZN(n802) );
  nd02d1 U578 ( .A1(n932), .A2(n802), .ZN(n866) );
  nd02d1 U582 ( .A1(n932), .A2(n931), .ZN(n807) );
  oai21d1 U583 ( .B1(n795), .B2(n807), .A(n806), .ZN(n808) );
  nd02d1 U586 ( .A1(n450), .A2(n429), .ZN(n814) );
  nr02d0 U587 ( .A1(n450), .A2(n429), .ZN(n815) );
  xr02d1 U595 ( .A1(n809), .A2(n867), .Z(product[12]) );
  nd02d1 U599 ( .A1(n928), .A2(n912), .ZN(n868) );
  oai21d1 U604 ( .B1(n809), .B2(n822), .A(n821), .ZN(n823) );
  nd02d1 U606 ( .A1(n500), .A2(n475), .ZN(n824) );
  nr02d0 U607 ( .A1(n500), .A2(n475), .ZN(n825) );
  nd02d1 U609 ( .A1(n753), .A2(n824), .ZN(n869) );
  oai21d1 U610 ( .B1(n821), .B2(n825), .A(n824), .ZN(n826) );
  nr02d0 U611 ( .A1(n822), .A2(n825), .ZN(n827) );
  xn02d1 U614 ( .A1(n823), .A2(n869), .ZN(product[14]) );
  nd02d1 U615 ( .A1(n528), .A2(n501), .ZN(n830) );
  nd02d1 U618 ( .A1(n927), .A2(n830), .ZN(n870) );
  xn02d1 U622 ( .A1(n829), .A2(n870), .ZN(product[15]) );
  nd02d1 U623 ( .A1(n556), .A2(n529), .ZN(n835) );
  nd02d1 U626 ( .A1(n929), .A2(n835), .ZN(n871) );
  nd02d1 U630 ( .A1(n929), .A2(n927), .ZN(n840) );
  oai21d1 U631 ( .B1(n828), .B2(n840), .A(n839), .ZN(n841) );
  invbd2 U650 ( .I(a[12]), .ZN(n44) );
  invbd2 U651 ( .I(b[1]), .ZN(n49) );
  ah01d0 U652 ( .A(n257), .B(n272), .CO(n453), .S(n452) );
  inv0d1 U653 ( .I(b[2]), .ZN(n50) );
  inv0d1 U654 ( .I(b[3]), .ZN(n51) );
  an02d1 U655 ( .A1(n474), .A2(n451), .Z(n908) );
  an02d1 U656 ( .A1(n924), .A2(n923), .Z(n909) );
  or02d1 U657 ( .A1(n65), .A2(n80), .Z(n910) );
  inv0d1 U658 ( .I(b[12]), .ZN(n911) );
  inv0d1 U659 ( .I(n908), .ZN(n912) );
  inv0d1 U660 ( .I(a[10]), .ZN(n913) );
  an02d1 U661 ( .A1(b[0]), .A2(a[13]), .Z(n272) );
  inv0d1 U662 ( .I(a[9]), .ZN(n41) );
  inv0d1 U663 ( .I(a[5]), .ZN(n37) );
  inv0d1 U664 ( .I(b[9]), .ZN(n57) );
  nd03d0 U665 ( .A1(n918), .A2(n919), .A3(n920), .ZN(n914) );
  nr02d0 U666 ( .A1(n51), .A2(n37), .ZN(n147) );
  inv0d1 U667 ( .I(a[2]), .ZN(n34) );
  inv0d1 U668 ( .I(b[5]), .ZN(n53) );
  nr02d0 U669 ( .A1(n53), .A2(n34), .ZN(n101) );
  inv0d1 U670 ( .I(a[8]), .ZN(n915) );
  ad01d0 U671 ( .A(n105), .B(n150), .CI(n135), .CO(n417), .S(n416) );
  inv0d1 U672 ( .I(b[11]), .ZN(n59) );
  inv0d1 U673 ( .I(a[6]), .ZN(n916) );
  nd02d1 U674 ( .A1(n922), .A2(n909), .ZN(n447) );
  ad01d0 U675 ( .A(n732), .B(n727), .CI(n851), .CO(n852), .S(product[27]) );
  ad01d0 U676 ( .A(n736), .B(n733), .CI(n852), .CO(n853), .S(product[28]) );
  nd02d0 U677 ( .A1(n412), .A2(n414), .ZN(n920) );
  ad01d0 U678 ( .A(n165), .B(n195), .CI(n180), .CO(n415), .S(n414) );
  inv0d1 U679 ( .I(b[6]), .ZN(n54) );
  xr02d1 U680 ( .A1(n414), .A2(n412), .Z(n917) );
  xr02d1 U681 ( .A1(n917), .A2(n416), .Z(n422) );
  nd02d0 U682 ( .A1(n416), .A2(n412), .ZN(n918) );
  nd02d1 U683 ( .A1(n416), .A2(n414), .ZN(n919) );
  nd03d0 U684 ( .A1(n918), .A2(n919), .A3(n920), .ZN(n423) );
  ad01d1 U685 ( .A(n75), .B(n210), .CI(n90), .CO(n413), .S(n412) );
  nd02d0 U686 ( .A1(n440), .A2(n914), .ZN(n922) );
  nr02d0 U687 ( .A1(n54), .A2(n38), .ZN(n166) );
  nr02d0 U688 ( .A1(n54), .A2(n36), .ZN(n134) );
  inv0d1 U689 ( .I(a[11]), .ZN(n43) );
  inv0d1 U690 ( .I(a[1]), .ZN(n33) );
  inv0d0 U691 ( .I(n828), .ZN(n829) );
  nd02d0 U692 ( .A1(n928), .A2(n813), .ZN(n822) );
  xr02d1 U693 ( .A1(n921), .A2(n868), .Z(product[13]) );
  ora21d1 U694 ( .B1(n809), .B2(n815), .A(n814), .Z(n921) );
  nd02d0 U695 ( .A1(n813), .A2(n814), .ZN(n867) );
  ad01d0 U696 ( .A(n430), .B(n413), .CI(n417), .CO(n441), .S(n440) );
  ad01d0 U697 ( .A(n395), .B(n399), .CI(n397), .CO(n421), .S(n420) );
  xr03d1 U698 ( .A1(n440), .A2(n421), .A3(n914), .Z(n446) );
  nd02d1 U699 ( .A1(n440), .A2(n421), .ZN(n923) );
  nd02d1 U700 ( .A1(n423), .A2(n421), .ZN(n924) );
  inv0d1 U701 ( .I(a[0]), .ZN(n925) );
  inv0d1 U702 ( .I(n830), .ZN(n832) );
  aoi21d1 U703 ( .B1(n808), .B2(n827), .A(n826), .ZN(n828) );
  inv0d1 U704 ( .I(n835), .ZN(n837) );
  xn02d1 U705 ( .A1(n926), .A2(n871), .ZN(product[16]) );
  aor21d1 U706 ( .B1(n829), .B2(n927), .A(n832), .Z(n926) );
  inv0d1 U707 ( .I(n825), .ZN(n753) );
  inv0d1 U708 ( .I(n808), .ZN(n809) );
  inv0d1 U709 ( .I(n795), .ZN(n796) );
  ad01d0 U710 ( .A(n583), .B(n606), .CI(n842), .CO(n843), .S(product[18]) );
  ad01d0 U711 ( .A(n607), .B(n628), .CI(n843), .CO(n844), .S(product[19]) );
  ad01d0 U712 ( .A(n629), .B(n648), .CI(n844), .CO(n845), .S(product[20]) );
  ad01d0 U713 ( .A(n557), .B(n582), .CI(n841), .CO(n842), .S(product[17]) );
  aoi21d1 U714 ( .B1(n929), .B2(n832), .A(n837), .ZN(n839) );
  aoi21d1 U715 ( .B1(n932), .B2(n799), .A(n804), .ZN(n806) );
  inv0d1 U716 ( .I(n802), .ZN(n804) );
  or02d1 U717 ( .A1(n528), .A2(n501), .Z(n927) );
  or02d1 U718 ( .A1(n474), .A2(n451), .Z(n928) );
  or02d1 U719 ( .A1(n556), .A2(n529), .Z(n929) );
  inv0d1 U720 ( .I(n815), .ZN(n813) );
  inv0d1 U721 ( .I(n797), .ZN(n799) );
  aoi21d1 U722 ( .B1(n786), .B2(n794), .A(n793), .ZN(n795) );
  aoi21d1 U723 ( .B1(n928), .B2(n812), .A(n908), .ZN(n821) );
  inv0d1 U724 ( .I(n814), .ZN(n812) );
  inv0d1 U725 ( .I(n792), .ZN(n748) );
  inv0d1 U726 ( .I(n789), .ZN(n747) );
  xn02d1 U727 ( .A1(n930), .A2(n866), .ZN(product[11]) );
  aor21d1 U728 ( .B1(n796), .B2(n931), .A(n799), .Z(n930) );
  inv0d1 U729 ( .I(n786), .ZN(n787) );
  inv0d1 U730 ( .I(n773), .ZN(n774) );
  ad01d0 U731 ( .A(n427), .B(n446), .CI(n448), .CO(n451), .S(n450) );
  ad01d0 U732 ( .A(n470), .B(n449), .CI(n472), .CO(n475), .S(n474) );
  ad01d0 U733 ( .A(n524), .B(n499), .CI(n526), .CO(n529), .S(n528) );
  ad01d0 U734 ( .A(n552), .B(n527), .CI(n554), .CO(n557), .S(n556) );
  ad01d0 U735 ( .A(n496), .B(n473), .CI(n498), .CO(n501), .S(n500) );
  ad01d0 U736 ( .A(n649), .B(n666), .CI(n845), .CO(n846), .S(product[21]) );
  ad01d0 U737 ( .A(n667), .B(n682), .CI(n846), .CO(n847), .S(product[22]) );
  ad01d0 U738 ( .A(n683), .B(n696), .CI(n847), .CO(n848), .S(product[23]) );
  ad01d0 U739 ( .A(n697), .B(n708), .CI(n848), .CO(n849), .S(product[24]) );
  ad01d0 U740 ( .A(n709), .B(n718), .CI(n849), .CO(n850), .S(product[25]) );
  ad01d0 U741 ( .A(n719), .B(n726), .CI(n850), .CO(n851), .S(product[26]) );
  aoi21d1 U742 ( .B1(n935), .B2(n777), .A(n782), .ZN(n784) );
  inv0d1 U743 ( .I(n780), .ZN(n782) );
  or02d1 U744 ( .A1(n408), .A2(n391), .Z(n931) );
  or02d1 U745 ( .A1(n428), .A2(n409), .Z(n932) );
  inv0d1 U746 ( .I(n775), .ZN(n777) );
  aoi21d1 U747 ( .B1(n768), .B2(n936), .A(n771), .ZN(n773) );
  inv0d1 U748 ( .I(n769), .ZN(n771) );
  ad01d0 U749 ( .A(n578), .B(n555), .CI(n580), .CO(n583), .S(n582) );
  ad01d0 U750 ( .A(n602), .B(n581), .CI(n604), .CO(n607), .S(n606) );
  ad01d0 U751 ( .A(n624), .B(n605), .CI(n626), .CO(n629), .S(n628) );
  ad01d0 U752 ( .A(n551), .B(n576), .CI(n553), .CO(n581), .S(n580) );
  ad01d0 U753 ( .A(n577), .B(n600), .CI(n579), .CO(n605), .S(n604) );
  ad01d0 U754 ( .A(n601), .B(n622), .CI(n603), .CO(n627), .S(n626) );
  ad01d0 U755 ( .A(n644), .B(n627), .CI(n646), .CO(n649), .S(n648) );
  xn02d1 U756 ( .A1(n933), .A2(n862), .ZN(product[7]) );
  aor21d1 U757 ( .B1(n774), .B2(n934), .A(n777), .Z(n933) );
  ad01d0 U758 ( .A(n514), .B(n491), .CI(n516), .CO(n523), .S(n522) );
  ad01d0 U759 ( .A(n488), .B(n490), .CI(n492), .CO(n497), .S(n496) );
  ad01d0 U760 ( .A(n521), .B(n546), .CI(n523), .CO(n553), .S(n552) );
  ad01d0 U761 ( .A(n443), .B(n464), .CI(n445), .CO(n471), .S(n470) );
  ad01d0 U762 ( .A(n493), .B(n518), .CI(n495), .CO(n525), .S(n524) );
  ad01d0 U763 ( .A(n404), .B(n389), .CI(n406), .CO(n409), .S(n408) );
  ad01d0 U764 ( .A(n424), .B(n407), .CI(n426), .CO(n429), .S(n428) );
  ad01d0 U765 ( .A(n359), .B(n370), .CI(n372), .CO(n375), .S(n374) );
  ad01d0 U766 ( .A(n347), .B(n356), .CI(n358), .CO(n361), .S(n360) );
  ad01d0 U767 ( .A(n373), .B(n386), .CI(n388), .CO(n391), .S(n390) );
  ad01d0 U768 ( .A(n400), .B(n387), .CI(n402), .CO(n407), .S(n406) );
  ad01d0 U769 ( .A(n442), .B(n444), .CI(n425), .CO(n449), .S(n448) );
  ad01d0 U770 ( .A(n420), .B(n405), .CI(n422), .CO(n427), .S(n426) );
  ad01d0 U771 ( .A(n519), .B(n542), .CI(n544), .CO(n551), .S(n550) );
  ad01d0 U772 ( .A(n466), .B(n447), .CI(n468), .CO(n473), .S(n472) );
  ad01d0 U773 ( .A(n469), .B(n471), .CI(n494), .CO(n499), .S(n498) );
  ad01d0 U774 ( .A(n548), .B(n525), .CI(n550), .CO(n555), .S(n554) );
  ad01d0 U775 ( .A(n520), .B(n522), .CI(n497), .CO(n527), .S(n526) );
  or02d1 U776 ( .A1(n348), .A2(n339), .Z(n934) );
  or02d1 U777 ( .A1(n360), .A2(n349), .Z(n935) );
  or02d1 U778 ( .A1(n338), .A2(n331), .Z(n936) );
  aoi21d1 U779 ( .B1(n937), .B2(n760), .A(n763), .ZN(n765) );
  inv0d1 U780 ( .I(n761), .ZN(n763) );
  ad01d0 U781 ( .A(n547), .B(n568), .CI(n570), .CO(n577), .S(n576) );
  ad01d0 U782 ( .A(n571), .B(n573), .CI(n594), .CO(n601), .S(n600) );
  ad01d0 U783 ( .A(n595), .B(n597), .CI(n616), .CO(n623), .S(n622) );
  ad01d0 U784 ( .A(n572), .B(n549), .CI(n574), .CO(n579), .S(n578) );
  ad01d0 U785 ( .A(n596), .B(n575), .CI(n598), .CO(n603), .S(n602) );
  ad01d0 U786 ( .A(n618), .B(n620), .CI(n599), .CO(n625), .S(n624) );
  ad01d0 U787 ( .A(n662), .B(n647), .CI(n664), .CO(n667), .S(n666) );
  ad01d0 U788 ( .A(n678), .B(n665), .CI(n680), .CO(n683), .S(n682) );
  ad01d0 U789 ( .A(n692), .B(n681), .CI(n694), .CO(n697), .S(n696) );
  ad01d0 U790 ( .A(n638), .B(n621), .CI(n640), .CO(n645), .S(n644) );
  ad01d0 U791 ( .A(n623), .B(n642), .CI(n625), .CO(n647), .S(n646) );
  ad01d0 U792 ( .A(n660), .B(n643), .CI(n645), .CO(n665), .S(n664) );
  ad01d0 U793 ( .A(n661), .B(n676), .CI(n663), .CO(n681), .S(n680) );
  ad01d0 U794 ( .A(n677), .B(n690), .CI(n679), .CO(n695), .S(n694) );
  ad01d0 U795 ( .A(n704), .B(n695), .CI(n706), .CO(n709), .S(n708) );
  ad01d0 U796 ( .A(n714), .B(n707), .CI(n716), .CO(n719), .S(n718) );
  ad01d0 U797 ( .A(n715), .B(n724), .CI(n717), .CO(n727), .S(n726) );
  inv0d1 U798 ( .I(n767), .ZN(n743) );
  inv0d1 U799 ( .I(n759), .ZN(n741) );
  ad01d0 U800 ( .A(n435), .B(n437), .CI(n460), .CO(n465), .S(n464) );
  ad01d0 U801 ( .A(n432), .B(n419), .CI(n438), .CO(n445), .S(n444) );
  ad01d0 U802 ( .A(n506), .B(n508), .CI(n504), .CO(n519), .S(n518) );
  ad01d0 U803 ( .A(n509), .B(n505), .CI(n511), .CO(n543), .S(n542) );
  ad01d0 U804 ( .A(n455), .B(n484), .CI(n482), .CO(n491), .S(n490) );
  ad01d0 U805 ( .A(n341), .B(n350), .CI(n343), .CO(n357), .S(n356) );
  ad01d0 U806 ( .A(n534), .B(n532), .CI(n513), .CO(n547), .S(n546) );
  ad01d0 U807 ( .A(n415), .B(n436), .CI(n434), .CO(n443), .S(n442) );
  ad01d0 U808 ( .A(n502), .B(n483), .CI(n479), .CO(n515), .S(n514) );
  ad01d0 U809 ( .A(n459), .B(n461), .CI(n457), .CO(n489), .S(n488) );
  ad01d0 U810 ( .A(n515), .B(n540), .CI(n517), .CO(n549), .S(n548) );
  ad01d0 U811 ( .A(n487), .B(n512), .CI(n489), .CO(n521), .S(n520) );
  ad01d0 U812 ( .A(n353), .B(n355), .CI(n366), .CO(n371), .S(n370) );
  ad01d0 U813 ( .A(n380), .B(n378), .CI(n369), .CO(n387), .S(n386) );
  ad01d0 U814 ( .A(n394), .B(n383), .CI(n385), .CO(n405), .S(n404) );
  ad01d0 U815 ( .A(n377), .B(n392), .CI(n379), .CO(n401), .S(n400) );
  ad01d0 U816 ( .A(n337), .B(n344), .CI(n346), .CO(n349), .S(n348) );
  ad01d0 U817 ( .A(n329), .B(n334), .CI(n336), .CO(n339), .S(n338) );
  ad01d0 U818 ( .A(n323), .B(n326), .CI(n328), .CO(n331), .S(n330) );
  ad01d0 U819 ( .A(n340), .B(n335), .CI(n342), .CO(n347), .S(n346) );
  ad01d0 U820 ( .A(n376), .B(n365), .CI(n367), .CO(n385), .S(n384) );
  ad01d0 U821 ( .A(n431), .B(n452), .CI(n433), .CO(n463), .S(n462) );
  ad01d0 U822 ( .A(n382), .B(n371), .CI(n384), .CO(n389), .S(n388) );
  ad01d0 U823 ( .A(n486), .B(n465), .CI(n467), .CO(n495), .S(n494) );
  ad01d0 U824 ( .A(n507), .B(n538), .CI(n536), .CO(n545), .S(n544) );
  ad01d0 U825 ( .A(n478), .B(n480), .CI(n463), .CO(n493), .S(n492) );
  ad01d0 U826 ( .A(n481), .B(n485), .CI(n510), .CO(n517), .S(n516) );
  ad01d0 U827 ( .A(n456), .B(n441), .CI(n462), .CO(n469), .S(n468) );
  ad01d0 U828 ( .A(n364), .B(n357), .CI(n368), .CO(n373), .S(n372) );
  ad01d0 U829 ( .A(n354), .B(n352), .CI(n345), .CO(n359), .S(n358) );
  ad01d0 U830 ( .A(n381), .B(n398), .CI(n396), .CO(n403), .S(n402) );
  ad01d0 U831 ( .A(n458), .B(n454), .CI(n439), .CO(n467), .S(n466) );
  ad01d0 U832 ( .A(n401), .B(n418), .CI(n403), .CO(n425), .S(n424) );
  ad01d0 U833 ( .A(n738), .B(n737), .CI(n853), .CO(n854), .S(product[29]) );
  or02d1 U834 ( .A1(n324), .A2(n322), .Z(n937) );
  ad01d0 U835 ( .A(n537), .B(n533), .CI(n539), .CO(n569), .S(n568) );
  ad01d0 U836 ( .A(n610), .B(n608), .CI(n593), .CO(n621), .S(n620) );
  ad01d0 U837 ( .A(n558), .B(n560), .CI(n541), .CO(n573), .S(n572) );
  ad01d0 U838 ( .A(n588), .B(n584), .CI(n567), .CO(n597), .S(n596) );
  ad01d0 U839 ( .A(n566), .B(n543), .CI(n545), .CO(n575), .S(n574) );
  ad01d0 U840 ( .A(n535), .B(n564), .CI(n562), .CO(n571), .S(n570) );
  ad01d0 U841 ( .A(n586), .B(n569), .CI(n592), .CO(n599), .S(n598) );
  ad01d0 U842 ( .A(n563), .B(n565), .CI(n590), .CO(n595), .S(n594) );
  ad01d0 U843 ( .A(n585), .B(n591), .CI(n589), .CO(n617), .S(n616) );
  ad01d0 U844 ( .A(n617), .B(n636), .CI(n619), .CO(n643), .S(n642) );
  ad01d0 U845 ( .A(n672), .B(n668), .CI(n670), .CO(n677), .S(n676) );
  ad01d0 U846 ( .A(n587), .B(n614), .CI(n612), .CO(n619), .S(n618) );
  ad01d0 U847 ( .A(n611), .B(n615), .CI(n613), .CO(n639), .S(n638) );
  ad01d0 U848 ( .A(n656), .B(n641), .CI(n658), .CO(n663), .S(n662) );
  ad01d0 U849 ( .A(n650), .B(n637), .CI(n639), .CO(n661), .S(n660) );
  ad01d0 U850 ( .A(n657), .B(n659), .CI(n674), .CO(n679), .S(n678) );
  ad01d0 U851 ( .A(n634), .B(n630), .CI(n632), .CO(n641), .S(n640) );
  ad01d0 U852 ( .A(n635), .B(n654), .CI(n652), .CO(n659), .S(n658) );
  ad01d0 U853 ( .A(n651), .B(n655), .CI(n653), .CO(n675), .S(n674) );
  ad01d0 U854 ( .A(n671), .B(n673), .CI(n686), .CO(n691), .S(n690) );
  ad01d0 U855 ( .A(n684), .B(n675), .CI(n688), .CO(n693), .S(n692) );
  ad01d0 U856 ( .A(n700), .B(n698), .CI(n689), .CO(n705), .S(n704) );
  ad01d0 U857 ( .A(n691), .B(n702), .CI(n693), .CO(n707), .S(n706) );
  ad01d0 U858 ( .A(n710), .B(n703), .CI(n705), .CO(n717), .S(n716) );
  ad01d0 U859 ( .A(n713), .B(n720), .CI(n722), .CO(n725), .S(n724) );
  ad01d0 U860 ( .A(n699), .B(n701), .CI(n712), .CO(n715), .S(n714) );
  ad01d0 U861 ( .A(n723), .B(n730), .CI(n725), .CO(n733), .S(n732) );
  ad01d0 U862 ( .A(n729), .B(n734), .CI(n731), .CO(n737), .S(n736) );
  an02d1 U863 ( .A1(n910), .A2(n756), .Z(product[1]) );
  ad01d0 U864 ( .A(n70), .B(n130), .CI(n85), .CO(n343), .S(n342) );
  ad01d0 U865 ( .A(n69), .B(n114), .CI(n99), .CO(n335), .S(n334) );
  ad01d0 U866 ( .A(n104), .B(n149), .CI(n119), .CO(n399), .S(n398) );
  ad01d0 U867 ( .A(n73), .B(n178), .CI(n88), .CO(n379), .S(n378) );
  ad01d0 U868 ( .A(n71), .B(n146), .CI(n86), .CO(n353), .S(n352) );
  ad01d0 U869 ( .A(n72), .B(n162), .CI(n87), .CO(n365), .S(n364) );
  ad01d0 U870 ( .A(n122), .B(n152), .CI(n137), .CO(n461), .S(n460) );
  ad01d0 U871 ( .A(n121), .B(n196), .CI(n181), .CO(n437), .S(n436) );
  ad01d0 U872 ( .A(n77), .B(n242), .CI(n92), .CO(n455), .S(n454) );
  ad01d0 U873 ( .A(n76), .B(n226), .CI(n211), .CO(n433), .S(n432) );
  ad01d0 U874 ( .A(n155), .B(n230), .CI(n185), .CO(n539), .S(n538) );
  ad01d0 U875 ( .A(n275), .B(n260), .CI(n245), .CO(n537), .S(n536) );
  ad01d0 U876 ( .A(n229), .B(n259), .CI(n244), .CO(n509), .S(n508) );
  ad01d0 U877 ( .A(n79), .B(n274), .CI(n94), .CO(n505), .S(n504) );
  ad01d0 U878 ( .A(n139), .B(n214), .CI(n184), .CO(n511), .S(n510) );
  ad01d0 U879 ( .A(n168), .B(n228), .CI(n93), .CO(n481), .S(n480) );
  ad01d0 U880 ( .A(n123), .B(n198), .CI(n153), .CO(n485), .S(n484) );
  ad01d0 U881 ( .A(n183), .B(n108), .CI(n213), .CO(n483), .S(n482) );
  ad01d0 U882 ( .A(n200), .B(n95), .CI(n110), .CO(n533), .S(n532) );
  ad01d0 U883 ( .A(n169), .B(n154), .CI(n477), .CO(n513), .S(n512) );
  ad01d0 U884 ( .A(n170), .B(n503), .CI(n530), .CO(n541), .S(n540) );
  ad01d0 U885 ( .A(n101), .B(n131), .CI(n116), .CO(n355), .S(n354) );
  ad01d0 U886 ( .A(n107), .B(n197), .CI(n167), .CO(n459), .S(n458) );
  ad01d0 U887 ( .A(n103), .B(n118), .CI(n363), .CO(n383), .S(n382) );
  ad01d0 U888 ( .A(n199), .B(n109), .CI(n124), .CO(n507), .S(n506) );
  ad01d0 U889 ( .A(n78), .B(n258), .CI(n243), .CO(n479), .S(n478) );
  ad01d0 U890 ( .A(n182), .B(n227), .CI(n212), .CO(n457), .S(n456) );
  ad01d0 U891 ( .A(n215), .B(n125), .CI(n140), .CO(n535), .S(n534) );
  ad01d0 U892 ( .A(n138), .B(n453), .CI(n476), .CO(n487), .S(n486) );
  ad01d0 U893 ( .A(n120), .B(n393), .CI(n410), .CO(n419), .S(n418) );
  ad01d0 U894 ( .A(n148), .B(n163), .CI(n133), .CO(n381), .S(n380) );
  ad01d0 U895 ( .A(n166), .B(n91), .CI(n106), .CO(n435), .S(n434) );
  ad01d0 U896 ( .A(n74), .B(n194), .CI(n179), .CO(n395), .S(n394) );
  ad01d0 U897 ( .A(n67), .B(n82), .CI(n321), .CO(n325), .S(n324) );
  ad01d0 U898 ( .A(n84), .B(n327), .CI(n332), .CO(n337), .S(n336) );
  ad01d0 U899 ( .A(n68), .B(n98), .CI(n83), .CO(n329), .S(n328) );
  ad01d0 U900 ( .A(n134), .B(n89), .CI(n164), .CO(n397), .S(n396) );
  ad01d0 U901 ( .A(n117), .B(n351), .CI(n362), .CO(n369), .S(n368) );
  ad01d0 U902 ( .A(n132), .B(n102), .CI(n147), .CO(n367), .S(n366) );
  ad01d0 U903 ( .A(n136), .B(n151), .CI(n411), .CO(n439), .S(n438) );
  ad01d0 U904 ( .A(n100), .B(n115), .CI(n333), .CO(n345), .S(n344) );
  ad01d0 U905 ( .A(n319), .B(n739), .CI(n854), .CO(product[31]), .S(
        product[30]) );
  ad01d0 U906 ( .A(n201), .B(n126), .CI(n276), .CO(n561), .S(n560) );
  ad01d0 U907 ( .A(n141), .B(n261), .CI(n156), .CO(n563), .S(n562) );
  ad01d0 U908 ( .A(n171), .B(n246), .CI(n231), .CO(n565), .S(n564) );
  ad01d0 U909 ( .A(n127), .B(n307), .CI(n142), .CO(n585), .S(n584) );
  ad01d0 U910 ( .A(n187), .B(n232), .CI(n217), .CO(n591), .S(n590) );
  ad01d0 U911 ( .A(n111), .B(n306), .CI(n291), .CO(n559), .S(n558) );
  ad01d0 U912 ( .A(n186), .B(n216), .CI(n531), .CO(n567), .S(n566) );
  ad01d0 U913 ( .A(n157), .B(n292), .CI(n277), .CO(n587), .S(n586) );
  ad01d0 U914 ( .A(n247), .B(n172), .CI(n262), .CO(n589), .S(n588) );
  ad01d0 U915 ( .A(n202), .B(n559), .CI(n561), .CO(n593), .S(n592) );
  ad01d0 U916 ( .A(n143), .B(n308), .CI(n293), .CO(n609), .S(n608) );
  ad01d0 U917 ( .A(n188), .B(n218), .CI(n203), .CO(n615), .S(n614) );
  ad01d0 U918 ( .A(n159), .B(n309), .CI(n294), .CO(n631), .S(n630) );
  ad01d0 U919 ( .A(n174), .B(n279), .CI(n264), .CO(n633), .S(n632) );
  ad01d0 U920 ( .A(n220), .B(n265), .CI(n250), .CO(n655), .S(n654) );
  ad01d0 U921 ( .A(n190), .B(n280), .CI(n205), .CO(n653), .S(n652) );
  ad01d0 U922 ( .A(n191), .B(n311), .CI(n296), .CO(n669), .S(n668) );
  ad01d0 U923 ( .A(n189), .B(n204), .CI(n609), .CO(n637), .S(n636) );
  ad01d0 U924 ( .A(n158), .B(n278), .CI(n263), .CO(n611), .S(n610) );
  ad01d0 U925 ( .A(n219), .B(n249), .CI(n234), .CO(n635), .S(n634) );
  ad01d0 U926 ( .A(n175), .B(n310), .CI(n295), .CO(n651), .S(n650) );
  ad01d0 U927 ( .A(n236), .B(n266), .CI(n251), .CO(n673), .S(n672) );
  ad01d0 U928 ( .A(n235), .B(n631), .CI(n633), .CO(n657), .S(n656) );
  ad01d0 U929 ( .A(n248), .B(n173), .CI(n233), .CO(n613), .S(n612) );
  ad01d0 U930 ( .A(n206), .B(n281), .CI(n221), .CO(n671), .S(n670) );
  ad01d0 U931 ( .A(n223), .B(n313), .CI(n298), .CO(n699), .S(n698) );
  ad01d0 U932 ( .A(n268), .B(n685), .CI(n687), .CO(n703), .S(n702) );
  ad01d0 U933 ( .A(n283), .B(n238), .CI(n253), .CO(n701), .S(n700) );
  ad01d0 U934 ( .A(n207), .B(n312), .CI(n297), .CO(n685), .S(n684) );
  ad01d0 U935 ( .A(n237), .B(n252), .CI(n669), .CO(n689), .S(n688) );
  ad01d0 U936 ( .A(n222), .B(n282), .CI(n267), .CO(n687), .S(n686) );
  ad01d0 U937 ( .A(n255), .B(n315), .CI(n300), .CO(n721), .S(n720) );
  ad01d0 U938 ( .A(n286), .B(n721), .CI(n728), .CO(n731), .S(n730) );
  ad01d0 U939 ( .A(n239), .B(n314), .CI(n299), .CO(n711), .S(n710) );
  ad01d0 U940 ( .A(n270), .B(n285), .CI(n711), .CO(n723), .S(n722) );
  ad01d0 U941 ( .A(n284), .B(n269), .CI(n254), .CO(n713), .S(n712) );
  ad01d0 U942 ( .A(n271), .B(n316), .CI(n301), .CO(n729), .S(n728) );
  ad01d0 U943 ( .A(n287), .B(n317), .CI(n302), .CO(n735), .S(n734) );
  ad01d0 U944 ( .A(n303), .B(n318), .CI(n735), .CO(n739), .S(n738) );
  inv0d1 U945 ( .I(a[0]), .ZN(n32) );
  inv0d1 U946 ( .I(a[3]), .ZN(n35) );
  inv0d1 U947 ( .I(a[4]), .ZN(n36) );
  inv0d1 U948 ( .I(a[6]), .ZN(n38) );
  inv0d1 U949 ( .I(a[7]), .ZN(n39) );
  inv0d1 U950 ( .I(a[8]), .ZN(n40) );
  inv0d1 U951 ( .I(a[10]), .ZN(n42) );
  inv0d1 U952 ( .I(a[13]), .ZN(n45) );
  inv0d1 U953 ( .I(a[14]), .ZN(n46) );
  inv0d1 U954 ( .I(a[15]), .ZN(n47) );
  inv0d1 U955 ( .I(b[0]), .ZN(n48) );
  inv0d1 U956 ( .I(b[4]), .ZN(n52) );
  inv0d1 U957 ( .I(b[7]), .ZN(n55) );
  inv0d1 U958 ( .I(b[8]), .ZN(n56) );
  inv0d1 U959 ( .I(b[10]), .ZN(n58) );
  inv0d1 U960 ( .I(b[12]), .ZN(n60) );
  inv0d1 U961 ( .I(b[13]), .ZN(n61) );
  inv0d1 U962 ( .I(b[14]), .ZN(n62) );
  inv0d1 U963 ( .I(b[15]), .ZN(n63) );
endmodule


module BLENDER_DW_mult_uns_5 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n741, n743, n747, n748, n753, n756, n758, n759, n760, n761, n763,
         n765, n766, n767, n768, n769, n771, n773, n774, n775, n777, n780,
         n782, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n799, n802, n804, n806, n807, n808, n809,
         n812, n813, n814, n815, n817, n819, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n832, n835, n837, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n908, n909, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933;

  nr02d0 U33 ( .A1(n48), .A2(n921), .ZN(product[0]) );
  nr02d0 U34 ( .A1(n49), .A2(n32), .ZN(n65) );
  nr02d0 U35 ( .A1(n50), .A2(n921), .ZN(n66) );
  nr02d0 U36 ( .A1(n51), .A2(n921), .ZN(n67) );
  nr02d0 U37 ( .A1(n52), .A2(n32), .ZN(n68) );
  nr02d0 U38 ( .A1(n53), .A2(n32), .ZN(n69) );
  nr02d0 U39 ( .A1(n54), .A2(n32), .ZN(n70) );
  nr02d0 U40 ( .A1(n55), .A2(n32), .ZN(n71) );
  nr02d0 U41 ( .A1(n56), .A2(n921), .ZN(n72) );
  nr02d0 U42 ( .A1(n57), .A2(n921), .ZN(n73) );
  nr02d0 U43 ( .A1(n58), .A2(n32), .ZN(n74) );
  nr02d0 U44 ( .A1(n59), .A2(n32), .ZN(n75) );
  nr02d0 U45 ( .A1(n60), .A2(n921), .ZN(n76) );
  nr02d0 U46 ( .A1(n61), .A2(n921), .ZN(n77) );
  nr02d0 U47 ( .A1(n62), .A2(n921), .ZN(n78) );
  nr02d0 U48 ( .A1(n63), .A2(n32), .ZN(n79) );
  nr02d0 U49 ( .A1(n48), .A2(n33), .ZN(n80) );
  nr02d0 U50 ( .A1(n49), .A2(n33), .ZN(n81) );
  nr02d0 U51 ( .A1(n50), .A2(n33), .ZN(n82) );
  nr02d0 U52 ( .A1(n51), .A2(n33), .ZN(n83) );
  nr02d0 U53 ( .A1(n52), .A2(n33), .ZN(n84) );
  nr02d0 U54 ( .A1(n53), .A2(n33), .ZN(n85) );
  nr02d0 U55 ( .A1(n54), .A2(n33), .ZN(n86) );
  nr02d0 U56 ( .A1(n55), .A2(n33), .ZN(n87) );
  nr02d0 U57 ( .A1(n56), .A2(n33), .ZN(n88) );
  nr02d0 U58 ( .A1(n57), .A2(n33), .ZN(n89) );
  nr02d0 U59 ( .A1(n58), .A2(n33), .ZN(n90) );
  nr02d0 U60 ( .A1(n59), .A2(n33), .ZN(n91) );
  nr02d0 U61 ( .A1(n60), .A2(n33), .ZN(n92) );
  nr02d0 U62 ( .A1(n61), .A2(n33), .ZN(n93) );
  nr02d0 U63 ( .A1(n62), .A2(n33), .ZN(n94) );
  nr02d0 U64 ( .A1(n63), .A2(n33), .ZN(n95) );
  nr02d0 U65 ( .A1(n48), .A2(n34), .ZN(n96) );
  nr02d0 U66 ( .A1(n49), .A2(n34), .ZN(n97) );
  nr02d0 U67 ( .A1(n50), .A2(n34), .ZN(n98) );
  nr02d0 U68 ( .A1(n51), .A2(n34), .ZN(n99) );
  nr02d0 U69 ( .A1(n52), .A2(n34), .ZN(n100) );
  nr02d0 U70 ( .A1(n53), .A2(n34), .ZN(n101) );
  nr02d0 U71 ( .A1(n54), .A2(n34), .ZN(n102) );
  nr02d0 U72 ( .A1(n55), .A2(n34), .ZN(n103) );
  nr02d0 U73 ( .A1(n56), .A2(n34), .ZN(n104) );
  nr02d0 U74 ( .A1(n57), .A2(n34), .ZN(n105) );
  nr02d0 U75 ( .A1(n58), .A2(n34), .ZN(n106) );
  nr02d0 U76 ( .A1(n59), .A2(n34), .ZN(n107) );
  nr02d0 U77 ( .A1(n60), .A2(n34), .ZN(n108) );
  nr02d0 U78 ( .A1(n61), .A2(n34), .ZN(n109) );
  nr02d0 U79 ( .A1(n62), .A2(n34), .ZN(n110) );
  nr02d0 U80 ( .A1(n63), .A2(n34), .ZN(n111) );
  nr02d0 U81 ( .A1(n48), .A2(n35), .ZN(n112) );
  nr02d0 U82 ( .A1(n49), .A2(n35), .ZN(n113) );
  nr02d0 U83 ( .A1(n50), .A2(n35), .ZN(n114) );
  nr02d0 U84 ( .A1(n51), .A2(n35), .ZN(n115) );
  nr02d0 U85 ( .A1(n52), .A2(n35), .ZN(n116) );
  nr02d0 U86 ( .A1(n53), .A2(n35), .ZN(n117) );
  nr02d0 U87 ( .A1(n54), .A2(n35), .ZN(n118) );
  nr02d0 U88 ( .A1(n55), .A2(n35), .ZN(n119) );
  nr02d0 U89 ( .A1(n56), .A2(n35), .ZN(n120) );
  nr02d0 U90 ( .A1(n57), .A2(n35), .ZN(n121) );
  nr02d0 U91 ( .A1(n58), .A2(n35), .ZN(n122) );
  nr02d0 U92 ( .A1(n59), .A2(n35), .ZN(n123) );
  nr02d0 U93 ( .A1(n60), .A2(n35), .ZN(n124) );
  nr02d0 U94 ( .A1(n61), .A2(n35), .ZN(n125) );
  nr02d0 U95 ( .A1(n62), .A2(n35), .ZN(n126) );
  nr02d0 U96 ( .A1(n63), .A2(n35), .ZN(n127) );
  nr02d0 U97 ( .A1(n48), .A2(n36), .ZN(n128) );
  nr02d0 U98 ( .A1(n49), .A2(n36), .ZN(n129) );
  nr02d0 U99 ( .A1(n50), .A2(n36), .ZN(n130) );
  nr02d0 U100 ( .A1(n51), .A2(n36), .ZN(n131) );
  nr02d0 U101 ( .A1(n52), .A2(n36), .ZN(n132) );
  nr02d0 U102 ( .A1(n53), .A2(n36), .ZN(n133) );
  nr02d0 U104 ( .A1(n55), .A2(n36), .ZN(n135) );
  nr02d0 U105 ( .A1(n56), .A2(n36), .ZN(n136) );
  nr02d0 U106 ( .A1(n57), .A2(n36), .ZN(n137) );
  nr02d0 U107 ( .A1(n58), .A2(n36), .ZN(n138) );
  nr02d0 U108 ( .A1(n59), .A2(n36), .ZN(n139) );
  nr02d0 U109 ( .A1(n60), .A2(n36), .ZN(n140) );
  nr02d0 U110 ( .A1(n61), .A2(n36), .ZN(n141) );
  nr02d0 U111 ( .A1(n62), .A2(n36), .ZN(n142) );
  nr02d0 U112 ( .A1(n63), .A2(n36), .ZN(n143) );
  nr02d0 U113 ( .A1(n48), .A2(n37), .ZN(n144) );
  nr02d0 U114 ( .A1(n49), .A2(n37), .ZN(n145) );
  nr02d0 U115 ( .A1(n50), .A2(n37), .ZN(n146) );
  nr02d0 U116 ( .A1(n51), .A2(n37), .ZN(n147) );
  nr02d0 U117 ( .A1(n52), .A2(n37), .ZN(n148) );
  nr02d0 U118 ( .A1(n53), .A2(n37), .ZN(n149) );
  nr02d0 U119 ( .A1(n54), .A2(n37), .ZN(n150) );
  nr02d0 U120 ( .A1(n55), .A2(n37), .ZN(n151) );
  nr02d0 U121 ( .A1(n56), .A2(n37), .ZN(n152) );
  nr02d0 U122 ( .A1(n57), .A2(n37), .ZN(n153) );
  nr02d0 U123 ( .A1(n58), .A2(n37), .ZN(n154) );
  nr02d0 U124 ( .A1(n59), .A2(n37), .ZN(n155) );
  nr02d0 U125 ( .A1(n60), .A2(n37), .ZN(n156) );
  nr02d0 U126 ( .A1(n61), .A2(n37), .ZN(n157) );
  nr02d0 U127 ( .A1(n62), .A2(n37), .ZN(n158) );
  nr02d0 U128 ( .A1(n63), .A2(n37), .ZN(n159) );
  nr02d0 U129 ( .A1(n48), .A2(n38), .ZN(n160) );
  nr02d0 U130 ( .A1(n49), .A2(n38), .ZN(n161) );
  nr02d0 U131 ( .A1(n50), .A2(n38), .ZN(n162) );
  nr02d0 U132 ( .A1(n51), .A2(n38), .ZN(n163) );
  nr02d0 U133 ( .A1(n52), .A2(n38), .ZN(n164) );
  nr02d0 U134 ( .A1(n53), .A2(n38), .ZN(n165) );
  nr02d0 U136 ( .A1(n55), .A2(n38), .ZN(n167) );
  nr02d0 U137 ( .A1(n56), .A2(n38), .ZN(n168) );
  nr02d0 U138 ( .A1(n57), .A2(n38), .ZN(n169) );
  nr02d0 U139 ( .A1(n58), .A2(n38), .ZN(n170) );
  nr02d0 U140 ( .A1(n59), .A2(n38), .ZN(n171) );
  nr02d0 U141 ( .A1(n60), .A2(n38), .ZN(n172) );
  nr02d0 U142 ( .A1(n61), .A2(n38), .ZN(n173) );
  nr02d0 U143 ( .A1(n62), .A2(n38), .ZN(n174) );
  nr02d0 U144 ( .A1(n63), .A2(n38), .ZN(n175) );
  nr02d0 U145 ( .A1(n48), .A2(n39), .ZN(n176) );
  nr02d0 U146 ( .A1(n49), .A2(n39), .ZN(n177) );
  nr02d0 U147 ( .A1(n50), .A2(n39), .ZN(n178) );
  nr02d0 U148 ( .A1(n51), .A2(n39), .ZN(n179) );
  nr02d0 U149 ( .A1(n52), .A2(n39), .ZN(n180) );
  nr02d0 U150 ( .A1(n53), .A2(n39), .ZN(n181) );
  nr02d0 U151 ( .A1(n54), .A2(n39), .ZN(n182) );
  nr02d0 U152 ( .A1(n55), .A2(n39), .ZN(n183) );
  nr02d0 U153 ( .A1(n56), .A2(n39), .ZN(n184) );
  nr02d0 U154 ( .A1(n57), .A2(n39), .ZN(n185) );
  nr02d0 U155 ( .A1(n58), .A2(n39), .ZN(n186) );
  nr02d0 U156 ( .A1(n59), .A2(n39), .ZN(n187) );
  nr02d0 U157 ( .A1(n60), .A2(n39), .ZN(n188) );
  nr02d0 U158 ( .A1(n61), .A2(n39), .ZN(n189) );
  nr02d0 U159 ( .A1(n62), .A2(n39), .ZN(n190) );
  nr02d0 U160 ( .A1(n63), .A2(n39), .ZN(n191) );
  nr02d0 U161 ( .A1(n48), .A2(n40), .ZN(n192) );
  nr02d0 U162 ( .A1(n49), .A2(n40), .ZN(n193) );
  nr02d0 U163 ( .A1(n50), .A2(n40), .ZN(n194) );
  nr02d0 U164 ( .A1(n51), .A2(n40), .ZN(n195) );
  nr02d0 U165 ( .A1(n52), .A2(n40), .ZN(n196) );
  nr02d0 U166 ( .A1(n53), .A2(n40), .ZN(n197) );
  nr02d0 U167 ( .A1(n54), .A2(n40), .ZN(n198) );
  nr02d0 U168 ( .A1(n55), .A2(n40), .ZN(n199) );
  nr02d0 U169 ( .A1(n56), .A2(n40), .ZN(n200) );
  nr02d0 U170 ( .A1(n57), .A2(n40), .ZN(n201) );
  nr02d0 U171 ( .A1(n58), .A2(n40), .ZN(n202) );
  nr02d0 U172 ( .A1(n59), .A2(n40), .ZN(n203) );
  nr02d0 U173 ( .A1(n60), .A2(n40), .ZN(n204) );
  nr02d0 U174 ( .A1(n61), .A2(n40), .ZN(n205) );
  nr02d0 U175 ( .A1(n62), .A2(n40), .ZN(n206) );
  nr02d0 U176 ( .A1(n63), .A2(n40), .ZN(n207) );
  nr02d0 U177 ( .A1(n48), .A2(n41), .ZN(n208) );
  nr02d0 U178 ( .A1(n49), .A2(n41), .ZN(n209) );
  nr02d0 U179 ( .A1(n50), .A2(n41), .ZN(n210) );
  nr02d0 U180 ( .A1(n51), .A2(n41), .ZN(n211) );
  nr02d0 U181 ( .A1(n52), .A2(n41), .ZN(n212) );
  nr02d0 U182 ( .A1(n53), .A2(n41), .ZN(n213) );
  nr02d0 U183 ( .A1(n54), .A2(n41), .ZN(n214) );
  nr02d0 U184 ( .A1(n55), .A2(n41), .ZN(n215) );
  nr02d0 U185 ( .A1(n56), .A2(n41), .ZN(n216) );
  nr02d0 U186 ( .A1(n57), .A2(n41), .ZN(n217) );
  nr02d0 U187 ( .A1(n58), .A2(n41), .ZN(n218) );
  nr02d0 U188 ( .A1(n59), .A2(n41), .ZN(n219) );
  nr02d0 U189 ( .A1(n60), .A2(n41), .ZN(n220) );
  nr02d0 U190 ( .A1(n61), .A2(n41), .ZN(n221) );
  nr02d0 U191 ( .A1(n62), .A2(n41), .ZN(n222) );
  nr02d0 U192 ( .A1(n63), .A2(n41), .ZN(n223) );
  nr02d0 U193 ( .A1(n48), .A2(n42), .ZN(n224) );
  nr02d0 U194 ( .A1(n49), .A2(n42), .ZN(n225) );
  nr02d0 U195 ( .A1(n50), .A2(n42), .ZN(n226) );
  nr02d0 U196 ( .A1(n51), .A2(n42), .ZN(n227) );
  nr02d0 U197 ( .A1(n52), .A2(n42), .ZN(n228) );
  nr02d0 U198 ( .A1(n53), .A2(n42), .ZN(n229) );
  nr02d0 U199 ( .A1(n54), .A2(n42), .ZN(n230) );
  nr02d0 U200 ( .A1(n55), .A2(n42), .ZN(n231) );
  nr02d0 U201 ( .A1(n56), .A2(n42), .ZN(n232) );
  nr02d0 U202 ( .A1(n57), .A2(n42), .ZN(n233) );
  nr02d0 U203 ( .A1(n58), .A2(n42), .ZN(n234) );
  nr02d0 U204 ( .A1(n59), .A2(n42), .ZN(n235) );
  nr02d0 U205 ( .A1(n60), .A2(n42), .ZN(n236) );
  nr02d0 U206 ( .A1(n61), .A2(n42), .ZN(n237) );
  nr02d0 U207 ( .A1(n62), .A2(n42), .ZN(n238) );
  nr02d0 U208 ( .A1(n63), .A2(n42), .ZN(n239) );
  nr02d0 U209 ( .A1(n48), .A2(n43), .ZN(n240) );
  nr02d0 U210 ( .A1(n49), .A2(n43), .ZN(n241) );
  nr02d0 U211 ( .A1(n50), .A2(n43), .ZN(n242) );
  nr02d0 U212 ( .A1(n51), .A2(n43), .ZN(n243) );
  nr02d0 U213 ( .A1(n52), .A2(n43), .ZN(n244) );
  nr02d0 U214 ( .A1(n53), .A2(n43), .ZN(n245) );
  nr02d0 U215 ( .A1(n54), .A2(n43), .ZN(n246) );
  nr02d0 U216 ( .A1(n55), .A2(n43), .ZN(n247) );
  nr02d0 U217 ( .A1(n56), .A2(n43), .ZN(n248) );
  nr02d0 U218 ( .A1(n57), .A2(n43), .ZN(n249) );
  nr02d0 U219 ( .A1(n58), .A2(n43), .ZN(n250) );
  nr02d0 U220 ( .A1(n59), .A2(n43), .ZN(n251) );
  nr02d0 U221 ( .A1(n60), .A2(n43), .ZN(n252) );
  nr02d0 U222 ( .A1(n61), .A2(n43), .ZN(n253) );
  nr02d0 U223 ( .A1(n62), .A2(n43), .ZN(n254) );
  nr02d0 U224 ( .A1(n63), .A2(n43), .ZN(n255) );
  nr02d0 U225 ( .A1(n48), .A2(n44), .ZN(n256) );
  nr02d0 U226 ( .A1(n49), .A2(n44), .ZN(n257) );
  nr02d0 U227 ( .A1(n50), .A2(n44), .ZN(n258) );
  nr02d0 U228 ( .A1(n51), .A2(n44), .ZN(n259) );
  nr02d0 U230 ( .A1(n53), .A2(n44), .ZN(n261) );
  nr02d0 U231 ( .A1(n54), .A2(n44), .ZN(n262) );
  nr02d0 U232 ( .A1(n55), .A2(n44), .ZN(n263) );
  nr02d0 U233 ( .A1(n56), .A2(n44), .ZN(n264) );
  nr02d0 U234 ( .A1(n57), .A2(n44), .ZN(n265) );
  nr02d0 U235 ( .A1(n58), .A2(n44), .ZN(n266) );
  nr02d0 U236 ( .A1(n59), .A2(n44), .ZN(n267) );
  nr02d0 U237 ( .A1(n60), .A2(n44), .ZN(n268) );
  nr02d0 U238 ( .A1(n61), .A2(n44), .ZN(n269) );
  nr02d0 U239 ( .A1(n62), .A2(n44), .ZN(n270) );
  nr02d0 U240 ( .A1(n63), .A2(n44), .ZN(n271) );
  nr02d0 U241 ( .A1(n48), .A2(n45), .ZN(n272) );
  nr02d0 U242 ( .A1(n49), .A2(n45), .ZN(n273) );
  nr02d0 U243 ( .A1(n50), .A2(n45), .ZN(n274) );
  nr02d0 U244 ( .A1(n51), .A2(n45), .ZN(n275) );
  nr02d0 U245 ( .A1(n52), .A2(n45), .ZN(n276) );
  nr02d0 U246 ( .A1(n53), .A2(n45), .ZN(n277) );
  nr02d0 U247 ( .A1(n54), .A2(n45), .ZN(n278) );
  nr02d0 U248 ( .A1(n55), .A2(n45), .ZN(n279) );
  nr02d0 U249 ( .A1(n56), .A2(n45), .ZN(n280) );
  nr02d0 U250 ( .A1(n57), .A2(n45), .ZN(n281) );
  nr02d0 U251 ( .A1(n58), .A2(n45), .ZN(n282) );
  nr02d0 U252 ( .A1(n59), .A2(n45), .ZN(n283) );
  nr02d0 U253 ( .A1(n60), .A2(n45), .ZN(n284) );
  nr02d0 U254 ( .A1(n61), .A2(n45), .ZN(n285) );
  nr02d0 U255 ( .A1(n62), .A2(n45), .ZN(n286) );
  nr02d0 U256 ( .A1(n63), .A2(n45), .ZN(n287) );
  nr02d0 U257 ( .A1(n48), .A2(n46), .ZN(n288) );
  nr02d0 U258 ( .A1(n49), .A2(n46), .ZN(n289) );
  nr02d0 U259 ( .A1(n50), .A2(n46), .ZN(n290) );
  nr02d0 U260 ( .A1(n51), .A2(n46), .ZN(n291) );
  nr02d0 U261 ( .A1(n52), .A2(n46), .ZN(n292) );
  nr02d0 U262 ( .A1(n53), .A2(n46), .ZN(n293) );
  nr02d0 U263 ( .A1(n54), .A2(n46), .ZN(n294) );
  nr02d0 U264 ( .A1(n55), .A2(n46), .ZN(n295) );
  nr02d0 U265 ( .A1(n56), .A2(n46), .ZN(n296) );
  nr02d0 U266 ( .A1(n57), .A2(n46), .ZN(n297) );
  nr02d0 U267 ( .A1(n58), .A2(n46), .ZN(n298) );
  nr02d0 U268 ( .A1(n59), .A2(n46), .ZN(n299) );
  nr02d0 U269 ( .A1(n60), .A2(n46), .ZN(n300) );
  nr02d0 U270 ( .A1(n61), .A2(n46), .ZN(n301) );
  nr02d0 U271 ( .A1(n62), .A2(n46), .ZN(n302) );
  nr02d0 U272 ( .A1(n63), .A2(n46), .ZN(n303) );
  nr02d0 U273 ( .A1(n48), .A2(n47), .ZN(n304) );
  nr02d0 U274 ( .A1(n49), .A2(n47), .ZN(n305) );
  nr02d0 U275 ( .A1(n50), .A2(n47), .ZN(n306) );
  nr02d0 U276 ( .A1(n51), .A2(n47), .ZN(n307) );
  nr02d0 U277 ( .A1(n52), .A2(n47), .ZN(n308) );
  nr02d0 U278 ( .A1(n53), .A2(n47), .ZN(n309) );
  nr02d0 U279 ( .A1(n54), .A2(n47), .ZN(n310) );
  nr02d0 U280 ( .A1(n55), .A2(n47), .ZN(n311) );
  nr02d0 U281 ( .A1(n56), .A2(n47), .ZN(n312) );
  nr02d0 U282 ( .A1(n57), .A2(n47), .ZN(n313) );
  nr02d0 U283 ( .A1(n58), .A2(n47), .ZN(n314) );
  nr02d0 U284 ( .A1(n59), .A2(n47), .ZN(n315) );
  nr02d0 U285 ( .A1(n60), .A2(n47), .ZN(n316) );
  nr02d0 U286 ( .A1(n61), .A2(n47), .ZN(n317) );
  nr02d0 U287 ( .A1(n62), .A2(n47), .ZN(n318) );
  nr02d0 U288 ( .A1(n63), .A2(n47), .ZN(n319) );
  ah01d0 U289 ( .A(n66), .B(n81), .CO(n321), .S(n320) );
  ah01d0 U290 ( .A(n97), .B(n112), .CO(n323), .S(n322) );
  ah01d0 U292 ( .A(n113), .B(n128), .CO(n327), .S(n326) );
  ah01d0 U295 ( .A(n129), .B(n144), .CO(n333), .S(n332) );
  ah01d0 U299 ( .A(n145), .B(n160), .CO(n341), .S(n340) );
  ah01d0 U304 ( .A(n161), .B(n176), .CO(n351), .S(n350) );
  ah01d0 U310 ( .A(n177), .B(n192), .CO(n363), .S(n362) );
  ah01d0 U317 ( .A(n193), .B(n208), .CO(n377), .S(n376) );
  ah01d0 U325 ( .A(n209), .B(n224), .CO(n393), .S(n392) );
  ah01d0 U334 ( .A(n225), .B(n240), .CO(n411), .S(n410) );
  ah01d0 U344 ( .A(n241), .B(n256), .CO(n431), .S(n430) );
  ah01d0 U367 ( .A(n273), .B(n288), .CO(n477), .S(n476) );
  ah01d0 U380 ( .A(n289), .B(n304), .CO(n503), .S(n502) );
  ah01d0 U394 ( .A(n290), .B(n305), .CO(n531), .S(n530) );
  nd02d1 U499 ( .A1(n65), .A2(n80), .ZN(n756) );
  nd02d1 U504 ( .A1(n320), .A2(n96), .ZN(n758) );
  nr02d0 U505 ( .A1(n320), .A2(n96), .ZN(n759) );
  nd02d1 U507 ( .A1(n741), .A2(n758), .ZN(n857) );
  oai21d1 U508 ( .B1(n759), .B2(n756), .A(n758), .ZN(n760) );
  xr02d1 U509 ( .A1(n857), .A2(n756), .Z(product[2]) );
  nd02d1 U510 ( .A1(n324), .A2(n322), .ZN(n761) );
  nd02d1 U513 ( .A1(n933), .A2(n761), .ZN(n858) );
  xn02d1 U517 ( .A1(n858), .A2(n760), .ZN(product[3]) );
  nd02d1 U518 ( .A1(n330), .A2(n325), .ZN(n766) );
  nr02d0 U519 ( .A1(n330), .A2(n325), .ZN(n767) );
  nd02d1 U521 ( .A1(n743), .A2(n766), .ZN(n859) );
  oai21d1 U522 ( .B1(n767), .B2(n765), .A(n766), .ZN(n768) );
  xr02d1 U523 ( .A1(n859), .A2(n765), .Z(product[4]) );
  nd02d1 U524 ( .A1(n338), .A2(n331), .ZN(n769) );
  nd02d1 U527 ( .A1(n932), .A2(n769), .ZN(n860) );
  xn02d1 U532 ( .A1(n860), .A2(n768), .ZN(product[5]) );
  nd02d1 U533 ( .A1(n348), .A2(n339), .ZN(n775) );
  nd02d1 U536 ( .A1(n930), .A2(n775), .ZN(n861) );
  xn02d1 U540 ( .A1(n861), .A2(n774), .ZN(product[6]) );
  nd02d1 U541 ( .A1(n360), .A2(n349), .ZN(n780) );
  nd02d1 U544 ( .A1(n931), .A2(n780), .ZN(n862) );
  nd02d1 U548 ( .A1(n931), .A2(n930), .ZN(n785) );
  oai21d1 U549 ( .B1(n785), .B2(n773), .A(n784), .ZN(n786) );
  nd02d1 U552 ( .A1(n374), .A2(n361), .ZN(n788) );
  nr02d0 U553 ( .A1(n374), .A2(n361), .ZN(n789) );
  nd02d1 U555 ( .A1(n747), .A2(n788), .ZN(n863) );
  oai21d1 U556 ( .B1(n787), .B2(n789), .A(n788), .ZN(n790) );
  xr02d1 U557 ( .A1(n787), .A2(n863), .Z(product[8]) );
  nd02d1 U558 ( .A1(n390), .A2(n375), .ZN(n791) );
  nr02d0 U559 ( .A1(n390), .A2(n375), .ZN(n792) );
  nd02d1 U561 ( .A1(n748), .A2(n791), .ZN(n864) );
  oai21d1 U562 ( .B1(n792), .B2(n788), .A(n791), .ZN(n793) );
  nr02d0 U563 ( .A1(n792), .A2(n789), .ZN(n794) );
  xn02d1 U566 ( .A1(n790), .A2(n864), .ZN(product[9]) );
  nd02d1 U567 ( .A1(n408), .A2(n391), .ZN(n797) );
  nd02d1 U570 ( .A1(n927), .A2(n797), .ZN(n865) );
  xn02d1 U574 ( .A1(n796), .A2(n865), .ZN(product[10]) );
  nd02d1 U575 ( .A1(n428), .A2(n409), .ZN(n802) );
  nd02d1 U578 ( .A1(n928), .A2(n802), .ZN(n866) );
  nd02d1 U582 ( .A1(n928), .A2(n927), .ZN(n807) );
  oai21d1 U583 ( .B1(n795), .B2(n807), .A(n806), .ZN(n808) );
  nd02d1 U586 ( .A1(n450), .A2(n429), .ZN(n814) );
  nr02d0 U587 ( .A1(n450), .A2(n429), .ZN(n815) );
  xr02d1 U595 ( .A1(n809), .A2(n867), .Z(product[12]) );
  nd02d1 U599 ( .A1(n924), .A2(n911), .ZN(n868) );
  oai21d1 U604 ( .B1(n809), .B2(n822), .A(n821), .ZN(n823) );
  nd02d1 U606 ( .A1(n500), .A2(n475), .ZN(n824) );
  nr02d0 U607 ( .A1(n500), .A2(n475), .ZN(n825) );
  nd02d1 U609 ( .A1(n753), .A2(n824), .ZN(n869) );
  oai21d1 U610 ( .B1(n821), .B2(n825), .A(n824), .ZN(n826) );
  nr02d0 U611 ( .A1(n822), .A2(n825), .ZN(n827) );
  xn02d1 U614 ( .A1(n823), .A2(n869), .ZN(product[14]) );
  nd02d1 U615 ( .A1(n528), .A2(n501), .ZN(n830) );
  nd02d1 U618 ( .A1(n923), .A2(n830), .ZN(n870) );
  xn02d1 U622 ( .A1(n829), .A2(n870), .ZN(product[15]) );
  nd02d1 U623 ( .A1(n556), .A2(n529), .ZN(n835) );
  nd02d1 U626 ( .A1(n925), .A2(n835), .ZN(n871) );
  nd02d1 U630 ( .A1(n925), .A2(n923), .ZN(n840) );
  oai21d1 U631 ( .B1(n828), .B2(n840), .A(n839), .ZN(n841) );
  ad01d1 U650 ( .A(n76), .B(n226), .CI(n211), .CO(n433), .S(n432) );
  ah01d1 U651 ( .A(n257), .B(n272), .CO(n453), .S(n452) );
  nr02d1 U652 ( .A1(n52), .A2(n44), .ZN(n260) );
  inv0d1 U653 ( .I(b[6]), .ZN(n54) );
  inv0d1 U654 ( .I(a[12]), .ZN(n44) );
  an02d1 U655 ( .A1(n920), .A2(n919), .Z(n908) );
  or02d1 U656 ( .A1(n65), .A2(n80), .Z(n909) );
  invbd2 U657 ( .I(n819), .ZN(n911) );
  ad01d0 U658 ( .A(n165), .B(n195), .CI(n180), .CO(n415), .S(n414) );
  inv0d1 U659 ( .I(b[2]), .ZN(n50) );
  nd02d0 U660 ( .A1(n474), .A2(n451), .ZN(n817) );
  inv0d1 U661 ( .I(a[2]), .ZN(n34) );
  ad01d0 U662 ( .A(n105), .B(n150), .CI(n135), .CO(n417), .S(n416) );
  inv0d1 U663 ( .I(a[9]), .ZN(n41) );
  inv0d1 U664 ( .I(a[5]), .ZN(n37) );
  inv0d1 U665 ( .I(b[9]), .ZN(n57) );
  inv0d1 U666 ( .I(b[11]), .ZN(n59) );
  nd03d0 U667 ( .A1(n914), .A2(n915), .A3(n916), .ZN(n912) );
  nd02d1 U668 ( .A1(n918), .A2(n908), .ZN(n447) );
  ad01d0 U669 ( .A(n732), .B(n727), .CI(n851), .CO(n852), .S(product[27]) );
  ad01d0 U670 ( .A(n736), .B(n733), .CI(n852), .CO(n853), .S(product[28]) );
  nd02d0 U671 ( .A1(n412), .A2(n414), .ZN(n916) );
  xr02d1 U672 ( .A1(n414), .A2(n412), .Z(n913) );
  xr02d1 U673 ( .A1(n913), .A2(n416), .Z(n422) );
  nd02d0 U674 ( .A1(n416), .A2(n412), .ZN(n914) );
  nd02d1 U675 ( .A1(n416), .A2(n414), .ZN(n915) );
  nd03d0 U676 ( .A1(n914), .A2(n915), .A3(n916), .ZN(n423) );
  ad01d1 U677 ( .A(n75), .B(n210), .CI(n90), .CO(n413), .S(n412) );
  nd02d0 U678 ( .A1(n440), .A2(n912), .ZN(n918) );
  nr02d0 U679 ( .A1(n54), .A2(n38), .ZN(n166) );
  nr02d0 U680 ( .A1(n54), .A2(n36), .ZN(n134) );
  inv0d1 U681 ( .I(a[11]), .ZN(n43) );
  inv0d1 U682 ( .I(a[1]), .ZN(n33) );
  inv0d0 U683 ( .I(n828), .ZN(n829) );
  nd02d0 U684 ( .A1(n924), .A2(n813), .ZN(n822) );
  xr02d1 U685 ( .A1(n917), .A2(n868), .Z(product[13]) );
  ora21d1 U686 ( .B1(n809), .B2(n815), .A(n814), .Z(n917) );
  nd02d0 U687 ( .A1(n813), .A2(n814), .ZN(n867) );
  ad01d0 U688 ( .A(n430), .B(n413), .CI(n417), .CO(n441), .S(n440) );
  ad01d0 U689 ( .A(n395), .B(n399), .CI(n397), .CO(n421), .S(n420) );
  xr03d1 U690 ( .A1(n440), .A2(n421), .A3(n912), .Z(n446) );
  nd02d1 U691 ( .A1(n440), .A2(n421), .ZN(n919) );
  nd02d1 U692 ( .A1(n423), .A2(n421), .ZN(n920) );
  inv0d1 U693 ( .I(a[0]), .ZN(n921) );
  inv0d1 U694 ( .I(n830), .ZN(n832) );
  aoi21d1 U695 ( .B1(n808), .B2(n827), .A(n826), .ZN(n828) );
  inv0d1 U696 ( .I(n835), .ZN(n837) );
  xn02d1 U697 ( .A1(n922), .A2(n871), .ZN(product[16]) );
  aor21d1 U698 ( .B1(n829), .B2(n923), .A(n832), .Z(n922) );
  inv0d1 U699 ( .I(n825), .ZN(n753) );
  inv0d1 U700 ( .I(n808), .ZN(n809) );
  inv0d1 U701 ( .I(n795), .ZN(n796) );
  ad01d0 U702 ( .A(n583), .B(n606), .CI(n842), .CO(n843), .S(product[18]) );
  ad01d0 U703 ( .A(n607), .B(n628), .CI(n843), .CO(n844), .S(product[19]) );
  ad01d0 U704 ( .A(n629), .B(n648), .CI(n844), .CO(n845), .S(product[20]) );
  ad01d0 U705 ( .A(n557), .B(n582), .CI(n841), .CO(n842), .S(product[17]) );
  aoi21d1 U706 ( .B1(n925), .B2(n832), .A(n837), .ZN(n839) );
  aoi21d1 U707 ( .B1(n928), .B2(n799), .A(n804), .ZN(n806) );
  inv0d1 U708 ( .I(n802), .ZN(n804) );
  or02d1 U709 ( .A1(n528), .A2(n501), .Z(n923) );
  or02d1 U710 ( .A1(n474), .A2(n451), .Z(n924) );
  or02d1 U711 ( .A1(n556), .A2(n529), .Z(n925) );
  inv0d1 U712 ( .I(n815), .ZN(n813) );
  inv0d1 U713 ( .I(n797), .ZN(n799) );
  aoi21d1 U714 ( .B1(n786), .B2(n794), .A(n793), .ZN(n795) );
  aoi21d1 U715 ( .B1(n924), .B2(n812), .A(n819), .ZN(n821) );
  inv0d1 U716 ( .I(n814), .ZN(n812) );
  inv0d1 U717 ( .I(n817), .ZN(n819) );
  inv0d1 U718 ( .I(n792), .ZN(n748) );
  inv0d1 U719 ( .I(n789), .ZN(n747) );
  xn02d1 U720 ( .A1(n926), .A2(n866), .ZN(product[11]) );
  aor21d1 U721 ( .B1(n796), .B2(n927), .A(n799), .Z(n926) );
  inv0d1 U722 ( .I(n786), .ZN(n787) );
  inv0d1 U723 ( .I(n773), .ZN(n774) );
  ad01d0 U724 ( .A(n427), .B(n446), .CI(n448), .CO(n451), .S(n450) );
  ad01d0 U725 ( .A(n470), .B(n449), .CI(n472), .CO(n475), .S(n474) );
  ad01d0 U726 ( .A(n524), .B(n499), .CI(n526), .CO(n529), .S(n528) );
  ad01d0 U727 ( .A(n552), .B(n527), .CI(n554), .CO(n557), .S(n556) );
  ad01d0 U728 ( .A(n496), .B(n473), .CI(n498), .CO(n501), .S(n500) );
  ad01d0 U729 ( .A(n649), .B(n666), .CI(n845), .CO(n846), .S(product[21]) );
  ad01d0 U730 ( .A(n667), .B(n682), .CI(n846), .CO(n847), .S(product[22]) );
  ad01d0 U731 ( .A(n683), .B(n696), .CI(n847), .CO(n848), .S(product[23]) );
  ad01d0 U732 ( .A(n697), .B(n708), .CI(n848), .CO(n849), .S(product[24]) );
  ad01d0 U733 ( .A(n709), .B(n718), .CI(n849), .CO(n850), .S(product[25]) );
  ad01d0 U734 ( .A(n719), .B(n726), .CI(n850), .CO(n851), .S(product[26]) );
  aoi21d1 U735 ( .B1(n931), .B2(n777), .A(n782), .ZN(n784) );
  inv0d1 U736 ( .I(n780), .ZN(n782) );
  or02d1 U737 ( .A1(n408), .A2(n391), .Z(n927) );
  or02d1 U738 ( .A1(n428), .A2(n409), .Z(n928) );
  inv0d1 U739 ( .I(n775), .ZN(n777) );
  aoi21d1 U740 ( .B1(n768), .B2(n932), .A(n771), .ZN(n773) );
  inv0d1 U741 ( .I(n769), .ZN(n771) );
  ad01d0 U742 ( .A(n578), .B(n555), .CI(n580), .CO(n583), .S(n582) );
  ad01d0 U743 ( .A(n602), .B(n581), .CI(n604), .CO(n607), .S(n606) );
  ad01d0 U744 ( .A(n624), .B(n605), .CI(n626), .CO(n629), .S(n628) );
  ad01d0 U745 ( .A(n551), .B(n576), .CI(n553), .CO(n581), .S(n580) );
  ad01d0 U746 ( .A(n577), .B(n600), .CI(n579), .CO(n605), .S(n604) );
  ad01d0 U747 ( .A(n601), .B(n622), .CI(n603), .CO(n627), .S(n626) );
  ad01d0 U748 ( .A(n644), .B(n627), .CI(n646), .CO(n649), .S(n648) );
  xn02d1 U749 ( .A1(n929), .A2(n862), .ZN(product[7]) );
  aor21d1 U750 ( .B1(n774), .B2(n930), .A(n777), .Z(n929) );
  ad01d0 U751 ( .A(n514), .B(n491), .CI(n516), .CO(n523), .S(n522) );
  ad01d0 U752 ( .A(n488), .B(n490), .CI(n492), .CO(n497), .S(n496) );
  ad01d0 U753 ( .A(n521), .B(n546), .CI(n523), .CO(n553), .S(n552) );
  ad01d0 U754 ( .A(n443), .B(n464), .CI(n445), .CO(n471), .S(n470) );
  ad01d0 U755 ( .A(n493), .B(n518), .CI(n495), .CO(n525), .S(n524) );
  ad01d0 U756 ( .A(n404), .B(n389), .CI(n406), .CO(n409), .S(n408) );
  ad01d0 U757 ( .A(n424), .B(n407), .CI(n426), .CO(n429), .S(n428) );
  ad01d0 U758 ( .A(n359), .B(n370), .CI(n372), .CO(n375), .S(n374) );
  ad01d0 U759 ( .A(n347), .B(n356), .CI(n358), .CO(n361), .S(n360) );
  ad01d0 U760 ( .A(n373), .B(n386), .CI(n388), .CO(n391), .S(n390) );
  ad01d0 U761 ( .A(n400), .B(n387), .CI(n402), .CO(n407), .S(n406) );
  ad01d0 U762 ( .A(n442), .B(n444), .CI(n425), .CO(n449), .S(n448) );
  ad01d0 U763 ( .A(n420), .B(n405), .CI(n422), .CO(n427), .S(n426) );
  ad01d0 U764 ( .A(n519), .B(n542), .CI(n544), .CO(n551), .S(n550) );
  ad01d0 U765 ( .A(n466), .B(n447), .CI(n468), .CO(n473), .S(n472) );
  ad01d0 U766 ( .A(n469), .B(n471), .CI(n494), .CO(n499), .S(n498) );
  ad01d0 U767 ( .A(n548), .B(n525), .CI(n550), .CO(n555), .S(n554) );
  ad01d0 U768 ( .A(n520), .B(n522), .CI(n497), .CO(n527), .S(n526) );
  or02d1 U769 ( .A1(n348), .A2(n339), .Z(n930) );
  or02d1 U770 ( .A1(n360), .A2(n349), .Z(n931) );
  or02d1 U771 ( .A1(n338), .A2(n331), .Z(n932) );
  aoi21d1 U772 ( .B1(n933), .B2(n760), .A(n763), .ZN(n765) );
  inv0d1 U773 ( .I(n761), .ZN(n763) );
  ad01d0 U774 ( .A(n547), .B(n568), .CI(n570), .CO(n577), .S(n576) );
  ad01d0 U775 ( .A(n571), .B(n573), .CI(n594), .CO(n601), .S(n600) );
  ad01d0 U776 ( .A(n595), .B(n597), .CI(n616), .CO(n623), .S(n622) );
  ad01d0 U777 ( .A(n572), .B(n549), .CI(n574), .CO(n579), .S(n578) );
  ad01d0 U778 ( .A(n596), .B(n575), .CI(n598), .CO(n603), .S(n602) );
  ad01d0 U779 ( .A(n618), .B(n620), .CI(n599), .CO(n625), .S(n624) );
  ad01d0 U780 ( .A(n662), .B(n647), .CI(n664), .CO(n667), .S(n666) );
  ad01d0 U781 ( .A(n678), .B(n665), .CI(n680), .CO(n683), .S(n682) );
  ad01d0 U782 ( .A(n692), .B(n681), .CI(n694), .CO(n697), .S(n696) );
  ad01d0 U783 ( .A(n638), .B(n621), .CI(n640), .CO(n645), .S(n644) );
  ad01d0 U784 ( .A(n623), .B(n642), .CI(n625), .CO(n647), .S(n646) );
  ad01d0 U785 ( .A(n660), .B(n643), .CI(n645), .CO(n665), .S(n664) );
  ad01d0 U786 ( .A(n661), .B(n676), .CI(n663), .CO(n681), .S(n680) );
  ad01d0 U787 ( .A(n677), .B(n690), .CI(n679), .CO(n695), .S(n694) );
  ad01d0 U788 ( .A(n704), .B(n695), .CI(n706), .CO(n709), .S(n708) );
  ad01d0 U789 ( .A(n714), .B(n707), .CI(n716), .CO(n719), .S(n718) );
  ad01d0 U790 ( .A(n715), .B(n724), .CI(n717), .CO(n727), .S(n726) );
  inv0d1 U791 ( .I(n767), .ZN(n743) );
  inv0d1 U792 ( .I(n759), .ZN(n741) );
  ad01d0 U793 ( .A(n435), .B(n437), .CI(n460), .CO(n465), .S(n464) );
  ad01d0 U794 ( .A(n432), .B(n419), .CI(n438), .CO(n445), .S(n444) );
  ad01d0 U795 ( .A(n506), .B(n508), .CI(n504), .CO(n519), .S(n518) );
  ad01d0 U796 ( .A(n509), .B(n505), .CI(n511), .CO(n543), .S(n542) );
  ad01d0 U797 ( .A(n455), .B(n484), .CI(n482), .CO(n491), .S(n490) );
  ad01d0 U798 ( .A(n341), .B(n350), .CI(n343), .CO(n357), .S(n356) );
  ad01d0 U799 ( .A(n534), .B(n532), .CI(n513), .CO(n547), .S(n546) );
  ad01d0 U800 ( .A(n415), .B(n436), .CI(n434), .CO(n443), .S(n442) );
  ad01d0 U801 ( .A(n502), .B(n483), .CI(n479), .CO(n515), .S(n514) );
  ad01d0 U802 ( .A(n459), .B(n461), .CI(n457), .CO(n489), .S(n488) );
  ad01d0 U803 ( .A(n515), .B(n540), .CI(n517), .CO(n549), .S(n548) );
  ad01d0 U804 ( .A(n487), .B(n512), .CI(n489), .CO(n521), .S(n520) );
  ad01d0 U805 ( .A(n353), .B(n355), .CI(n366), .CO(n371), .S(n370) );
  ad01d0 U806 ( .A(n380), .B(n378), .CI(n369), .CO(n387), .S(n386) );
  ad01d0 U807 ( .A(n394), .B(n383), .CI(n385), .CO(n405), .S(n404) );
  ad01d0 U808 ( .A(n377), .B(n392), .CI(n379), .CO(n401), .S(n400) );
  ad01d0 U809 ( .A(n337), .B(n344), .CI(n346), .CO(n349), .S(n348) );
  ad01d0 U810 ( .A(n329), .B(n334), .CI(n336), .CO(n339), .S(n338) );
  ad01d0 U811 ( .A(n323), .B(n326), .CI(n328), .CO(n331), .S(n330) );
  ad01d0 U812 ( .A(n340), .B(n335), .CI(n342), .CO(n347), .S(n346) );
  ad01d0 U813 ( .A(n376), .B(n365), .CI(n367), .CO(n385), .S(n384) );
  ad01d0 U814 ( .A(n431), .B(n452), .CI(n433), .CO(n463), .S(n462) );
  ad01d0 U815 ( .A(n382), .B(n371), .CI(n384), .CO(n389), .S(n388) );
  ad01d0 U816 ( .A(n486), .B(n465), .CI(n467), .CO(n495), .S(n494) );
  ad01d0 U817 ( .A(n507), .B(n538), .CI(n536), .CO(n545), .S(n544) );
  ad01d0 U818 ( .A(n478), .B(n480), .CI(n463), .CO(n493), .S(n492) );
  ad01d0 U819 ( .A(n481), .B(n485), .CI(n510), .CO(n517), .S(n516) );
  ad01d0 U820 ( .A(n456), .B(n441), .CI(n462), .CO(n469), .S(n468) );
  ad01d0 U821 ( .A(n364), .B(n357), .CI(n368), .CO(n373), .S(n372) );
  ad01d0 U822 ( .A(n354), .B(n352), .CI(n345), .CO(n359), .S(n358) );
  ad01d0 U823 ( .A(n381), .B(n398), .CI(n396), .CO(n403), .S(n402) );
  ad01d0 U824 ( .A(n458), .B(n454), .CI(n439), .CO(n467), .S(n466) );
  ad01d0 U825 ( .A(n401), .B(n418), .CI(n403), .CO(n425), .S(n424) );
  ad01d0 U826 ( .A(n738), .B(n737), .CI(n853), .CO(n854), .S(product[29]) );
  or02d1 U827 ( .A1(n324), .A2(n322), .Z(n933) );
  ad01d0 U828 ( .A(n537), .B(n533), .CI(n539), .CO(n569), .S(n568) );
  ad01d0 U829 ( .A(n610), .B(n608), .CI(n593), .CO(n621), .S(n620) );
  ad01d0 U830 ( .A(n558), .B(n560), .CI(n541), .CO(n573), .S(n572) );
  ad01d0 U831 ( .A(n588), .B(n584), .CI(n567), .CO(n597), .S(n596) );
  ad01d0 U832 ( .A(n566), .B(n543), .CI(n545), .CO(n575), .S(n574) );
  ad01d0 U833 ( .A(n535), .B(n564), .CI(n562), .CO(n571), .S(n570) );
  ad01d0 U834 ( .A(n586), .B(n569), .CI(n592), .CO(n599), .S(n598) );
  ad01d0 U835 ( .A(n563), .B(n565), .CI(n590), .CO(n595), .S(n594) );
  ad01d0 U836 ( .A(n585), .B(n591), .CI(n589), .CO(n617), .S(n616) );
  ad01d0 U837 ( .A(n617), .B(n636), .CI(n619), .CO(n643), .S(n642) );
  ad01d0 U838 ( .A(n672), .B(n668), .CI(n670), .CO(n677), .S(n676) );
  ad01d0 U839 ( .A(n587), .B(n614), .CI(n612), .CO(n619), .S(n618) );
  ad01d0 U840 ( .A(n611), .B(n615), .CI(n613), .CO(n639), .S(n638) );
  ad01d0 U841 ( .A(n656), .B(n641), .CI(n658), .CO(n663), .S(n662) );
  ad01d0 U842 ( .A(n650), .B(n637), .CI(n639), .CO(n661), .S(n660) );
  ad01d0 U843 ( .A(n657), .B(n659), .CI(n674), .CO(n679), .S(n678) );
  ad01d0 U844 ( .A(n634), .B(n630), .CI(n632), .CO(n641), .S(n640) );
  ad01d0 U845 ( .A(n635), .B(n654), .CI(n652), .CO(n659), .S(n658) );
  ad01d0 U846 ( .A(n651), .B(n655), .CI(n653), .CO(n675), .S(n674) );
  ad01d0 U847 ( .A(n671), .B(n673), .CI(n686), .CO(n691), .S(n690) );
  ad01d0 U848 ( .A(n684), .B(n675), .CI(n688), .CO(n693), .S(n692) );
  ad01d0 U849 ( .A(n700), .B(n698), .CI(n689), .CO(n705), .S(n704) );
  ad01d0 U850 ( .A(n691), .B(n702), .CI(n693), .CO(n707), .S(n706) );
  ad01d0 U851 ( .A(n710), .B(n703), .CI(n705), .CO(n717), .S(n716) );
  ad01d0 U852 ( .A(n713), .B(n720), .CI(n722), .CO(n725), .S(n724) );
  ad01d0 U853 ( .A(n699), .B(n701), .CI(n712), .CO(n715), .S(n714) );
  ad01d0 U854 ( .A(n723), .B(n730), .CI(n725), .CO(n733), .S(n732) );
  ad01d0 U855 ( .A(n729), .B(n734), .CI(n731), .CO(n737), .S(n736) );
  an02d1 U856 ( .A1(n909), .A2(n756), .Z(product[1]) );
  ad01d0 U857 ( .A(n70), .B(n130), .CI(n85), .CO(n343), .S(n342) );
  ad01d0 U858 ( .A(n69), .B(n114), .CI(n99), .CO(n335), .S(n334) );
  ad01d0 U859 ( .A(n104), .B(n149), .CI(n119), .CO(n399), .S(n398) );
  ad01d0 U860 ( .A(n73), .B(n178), .CI(n88), .CO(n379), .S(n378) );
  ad01d0 U861 ( .A(n71), .B(n146), .CI(n86), .CO(n353), .S(n352) );
  ad01d0 U862 ( .A(n72), .B(n162), .CI(n87), .CO(n365), .S(n364) );
  ad01d0 U863 ( .A(n122), .B(n152), .CI(n137), .CO(n461), .S(n460) );
  ad01d0 U864 ( .A(n121), .B(n196), .CI(n181), .CO(n437), .S(n436) );
  ad01d0 U865 ( .A(n77), .B(n242), .CI(n92), .CO(n455), .S(n454) );
  ad01d0 U866 ( .A(n155), .B(n230), .CI(n185), .CO(n539), .S(n538) );
  ad01d0 U867 ( .A(n275), .B(n260), .CI(n245), .CO(n537), .S(n536) );
  ad01d0 U868 ( .A(n229), .B(n259), .CI(n244), .CO(n509), .S(n508) );
  ad01d0 U869 ( .A(n79), .B(n274), .CI(n94), .CO(n505), .S(n504) );
  ad01d0 U870 ( .A(n139), .B(n214), .CI(n184), .CO(n511), .S(n510) );
  ad01d0 U871 ( .A(n168), .B(n228), .CI(n93), .CO(n481), .S(n480) );
  ad01d0 U872 ( .A(n123), .B(n198), .CI(n153), .CO(n485), .S(n484) );
  ad01d0 U873 ( .A(n183), .B(n108), .CI(n213), .CO(n483), .S(n482) );
  ad01d0 U874 ( .A(n200), .B(n95), .CI(n110), .CO(n533), .S(n532) );
  ad01d0 U875 ( .A(n169), .B(n154), .CI(n477), .CO(n513), .S(n512) );
  ad01d0 U876 ( .A(n170), .B(n503), .CI(n530), .CO(n541), .S(n540) );
  ad01d0 U877 ( .A(n101), .B(n131), .CI(n116), .CO(n355), .S(n354) );
  ad01d0 U878 ( .A(n107), .B(n197), .CI(n167), .CO(n459), .S(n458) );
  ad01d0 U879 ( .A(n103), .B(n118), .CI(n363), .CO(n383), .S(n382) );
  ad01d0 U880 ( .A(n199), .B(n109), .CI(n124), .CO(n507), .S(n506) );
  ad01d0 U881 ( .A(n78), .B(n258), .CI(n243), .CO(n479), .S(n478) );
  ad01d0 U882 ( .A(n182), .B(n227), .CI(n212), .CO(n457), .S(n456) );
  ad01d0 U883 ( .A(n215), .B(n125), .CI(n140), .CO(n535), .S(n534) );
  ad01d0 U884 ( .A(n138), .B(n453), .CI(n476), .CO(n487), .S(n486) );
  ad01d0 U885 ( .A(n120), .B(n393), .CI(n410), .CO(n419), .S(n418) );
  ad01d0 U886 ( .A(n148), .B(n163), .CI(n133), .CO(n381), .S(n380) );
  ad01d0 U887 ( .A(n166), .B(n91), .CI(n106), .CO(n435), .S(n434) );
  ad01d0 U888 ( .A(n74), .B(n194), .CI(n179), .CO(n395), .S(n394) );
  ad01d0 U889 ( .A(n67), .B(n82), .CI(n321), .CO(n325), .S(n324) );
  ad01d0 U890 ( .A(n84), .B(n327), .CI(n332), .CO(n337), .S(n336) );
  ad01d0 U891 ( .A(n68), .B(n98), .CI(n83), .CO(n329), .S(n328) );
  ad01d0 U892 ( .A(n134), .B(n89), .CI(n164), .CO(n397), .S(n396) );
  ad01d0 U893 ( .A(n117), .B(n351), .CI(n362), .CO(n369), .S(n368) );
  ad01d0 U894 ( .A(n132), .B(n102), .CI(n147), .CO(n367), .S(n366) );
  ad01d0 U895 ( .A(n136), .B(n151), .CI(n411), .CO(n439), .S(n438) );
  ad01d0 U896 ( .A(n100), .B(n115), .CI(n333), .CO(n345), .S(n344) );
  ad01d0 U897 ( .A(n319), .B(n739), .CI(n854), .CO(product[31]), .S(
        product[30]) );
  ad01d0 U898 ( .A(n201), .B(n126), .CI(n276), .CO(n561), .S(n560) );
  ad01d0 U899 ( .A(n141), .B(n261), .CI(n156), .CO(n563), .S(n562) );
  ad01d0 U900 ( .A(n171), .B(n246), .CI(n231), .CO(n565), .S(n564) );
  ad01d0 U901 ( .A(n127), .B(n307), .CI(n142), .CO(n585), .S(n584) );
  ad01d0 U902 ( .A(n187), .B(n232), .CI(n217), .CO(n591), .S(n590) );
  ad01d0 U903 ( .A(n111), .B(n306), .CI(n291), .CO(n559), .S(n558) );
  ad01d0 U904 ( .A(n186), .B(n216), .CI(n531), .CO(n567), .S(n566) );
  ad01d0 U905 ( .A(n157), .B(n292), .CI(n277), .CO(n587), .S(n586) );
  ad01d0 U906 ( .A(n247), .B(n172), .CI(n262), .CO(n589), .S(n588) );
  ad01d0 U907 ( .A(n202), .B(n559), .CI(n561), .CO(n593), .S(n592) );
  ad01d0 U908 ( .A(n143), .B(n308), .CI(n293), .CO(n609), .S(n608) );
  ad01d0 U909 ( .A(n188), .B(n218), .CI(n203), .CO(n615), .S(n614) );
  ad01d0 U910 ( .A(n159), .B(n309), .CI(n294), .CO(n631), .S(n630) );
  ad01d0 U911 ( .A(n174), .B(n279), .CI(n264), .CO(n633), .S(n632) );
  ad01d0 U912 ( .A(n220), .B(n265), .CI(n250), .CO(n655), .S(n654) );
  ad01d0 U913 ( .A(n190), .B(n280), .CI(n205), .CO(n653), .S(n652) );
  ad01d0 U914 ( .A(n191), .B(n311), .CI(n296), .CO(n669), .S(n668) );
  ad01d0 U915 ( .A(n189), .B(n204), .CI(n609), .CO(n637), .S(n636) );
  ad01d0 U916 ( .A(n158), .B(n278), .CI(n263), .CO(n611), .S(n610) );
  ad01d0 U917 ( .A(n219), .B(n249), .CI(n234), .CO(n635), .S(n634) );
  ad01d0 U918 ( .A(n175), .B(n310), .CI(n295), .CO(n651), .S(n650) );
  ad01d0 U919 ( .A(n236), .B(n266), .CI(n251), .CO(n673), .S(n672) );
  ad01d0 U920 ( .A(n235), .B(n631), .CI(n633), .CO(n657), .S(n656) );
  ad01d0 U921 ( .A(n248), .B(n173), .CI(n233), .CO(n613), .S(n612) );
  ad01d0 U922 ( .A(n206), .B(n281), .CI(n221), .CO(n671), .S(n670) );
  ad01d0 U923 ( .A(n223), .B(n313), .CI(n298), .CO(n699), .S(n698) );
  ad01d0 U924 ( .A(n268), .B(n685), .CI(n687), .CO(n703), .S(n702) );
  ad01d0 U925 ( .A(n283), .B(n238), .CI(n253), .CO(n701), .S(n700) );
  ad01d0 U926 ( .A(n207), .B(n312), .CI(n297), .CO(n685), .S(n684) );
  ad01d0 U927 ( .A(n237), .B(n252), .CI(n669), .CO(n689), .S(n688) );
  ad01d0 U928 ( .A(n222), .B(n282), .CI(n267), .CO(n687), .S(n686) );
  ad01d0 U929 ( .A(n255), .B(n315), .CI(n300), .CO(n721), .S(n720) );
  ad01d0 U930 ( .A(n286), .B(n721), .CI(n728), .CO(n731), .S(n730) );
  ad01d0 U931 ( .A(n239), .B(n314), .CI(n299), .CO(n711), .S(n710) );
  ad01d0 U932 ( .A(n270), .B(n285), .CI(n711), .CO(n723), .S(n722) );
  ad01d0 U933 ( .A(n284), .B(n269), .CI(n254), .CO(n713), .S(n712) );
  ad01d0 U934 ( .A(n271), .B(n316), .CI(n301), .CO(n729), .S(n728) );
  ad01d0 U935 ( .A(n287), .B(n317), .CI(n302), .CO(n735), .S(n734) );
  ad01d0 U936 ( .A(n303), .B(n318), .CI(n735), .CO(n739), .S(n738) );
  inv0d1 U937 ( .I(a[0]), .ZN(n32) );
  inv0d1 U938 ( .I(a[3]), .ZN(n35) );
  inv0d1 U939 ( .I(a[4]), .ZN(n36) );
  inv0d1 U940 ( .I(a[6]), .ZN(n38) );
  inv0d1 U941 ( .I(a[7]), .ZN(n39) );
  inv0d1 U942 ( .I(a[8]), .ZN(n40) );
  inv0d1 U943 ( .I(a[10]), .ZN(n42) );
  inv0d1 U944 ( .I(a[13]), .ZN(n45) );
  inv0d1 U945 ( .I(a[14]), .ZN(n46) );
  inv0d1 U946 ( .I(a[15]), .ZN(n47) );
  inv0d1 U947 ( .I(b[0]), .ZN(n48) );
  inv0d1 U948 ( .I(b[1]), .ZN(n49) );
  inv0d1 U949 ( .I(b[3]), .ZN(n51) );
  inv0d1 U950 ( .I(b[4]), .ZN(n52) );
  inv0d1 U951 ( .I(b[5]), .ZN(n53) );
  inv0d1 U952 ( .I(b[7]), .ZN(n55) );
  inv0d1 U953 ( .I(b[8]), .ZN(n56) );
  inv0d1 U954 ( .I(b[10]), .ZN(n58) );
  inv0d1 U955 ( .I(b[12]), .ZN(n60) );
  inv0d1 U956 ( .I(b[13]), .ZN(n61) );
  inv0d1 U957 ( .I(b[14]), .ZN(n62) );
  inv0d1 U958 ( .I(b[15]), .ZN(n63) );
endmodule


module BLENDER_DW_mult_uns_3 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432;

  nr02d0 U25 ( .A1(n36), .A2(n24), .ZN(product[0]) );
  nr02d0 U26 ( .A1(n37), .A2(n24), .ZN(n49) );
  nr02d0 U27 ( .A1(n38), .A2(n24), .ZN(n50) );
  nr02d0 U28 ( .A1(n39), .A2(n24), .ZN(n51) );
  nr02d0 U29 ( .A1(n40), .A2(n24), .ZN(n52) );
  nr02d0 U30 ( .A1(n41), .A2(n24), .ZN(n53) );
  nr02d0 U31 ( .A1(n42), .A2(n24), .ZN(n54) );
  nr02d0 U32 ( .A1(n43), .A2(n24), .ZN(n55) );
  nr02d0 U33 ( .A1(n44), .A2(n24), .ZN(n56) );
  nr02d0 U34 ( .A1(n45), .A2(n24), .ZN(n57) );
  nr02d0 U35 ( .A1(n46), .A2(n24), .ZN(n58) );
  nr02d0 U36 ( .A1(n47), .A2(n24), .ZN(n59) );
  nr02d0 U37 ( .A1(n36), .A2(n25), .ZN(n60) );
  nr02d0 U38 ( .A1(n37), .A2(n25), .ZN(n61) );
  nr02d0 U39 ( .A1(n38), .A2(n25), .ZN(n62) );
  nr02d0 U40 ( .A1(n39), .A2(n25), .ZN(n63) );
  nr02d0 U41 ( .A1(n40), .A2(n25), .ZN(n64) );
  nr02d0 U42 ( .A1(n41), .A2(n25), .ZN(n65) );
  nr02d0 U43 ( .A1(n42), .A2(n25), .ZN(n66) );
  nr02d0 U44 ( .A1(n43), .A2(n25), .ZN(n67) );
  nr02d0 U45 ( .A1(n44), .A2(n25), .ZN(n68) );
  nr02d0 U46 ( .A1(n45), .A2(n25), .ZN(n69) );
  nr02d0 U47 ( .A1(n46), .A2(n25), .ZN(n70) );
  nr02d0 U48 ( .A1(n47), .A2(n25), .ZN(n71) );
  nr02d0 U49 ( .A1(n36), .A2(n26), .ZN(n72) );
  nr02d0 U50 ( .A1(n37), .A2(n26), .ZN(n73) );
  nr02d0 U51 ( .A1(n38), .A2(n26), .ZN(n74) );
  nr02d0 U52 ( .A1(n39), .A2(n26), .ZN(n75) );
  nr02d0 U53 ( .A1(n40), .A2(n26), .ZN(n76) );
  nr02d0 U54 ( .A1(n41), .A2(n26), .ZN(n77) );
  nr02d0 U55 ( .A1(n42), .A2(n26), .ZN(n78) );
  nr02d0 U56 ( .A1(n43), .A2(n26), .ZN(n79) );
  nr02d0 U57 ( .A1(n44), .A2(n26), .ZN(n80) );
  nr02d0 U58 ( .A1(n45), .A2(n26), .ZN(n81) );
  nr02d0 U59 ( .A1(n46), .A2(n26), .ZN(n82) );
  nr02d0 U60 ( .A1(n47), .A2(n26), .ZN(n83) );
  nr02d0 U61 ( .A1(n36), .A2(n27), .ZN(n84) );
  nr02d0 U62 ( .A1(n37), .A2(n27), .ZN(n85) );
  nr02d0 U63 ( .A1(n38), .A2(n27), .ZN(n86) );
  nr02d0 U64 ( .A1(n39), .A2(n27), .ZN(n87) );
  nr02d0 U65 ( .A1(n40), .A2(n27), .ZN(n88) );
  nr02d0 U66 ( .A1(n41), .A2(n27), .ZN(n89) );
  nr02d0 U67 ( .A1(n42), .A2(n27), .ZN(n90) );
  nr02d0 U68 ( .A1(n43), .A2(n27), .ZN(n91) );
  nr02d0 U69 ( .A1(n44), .A2(n27), .ZN(n92) );
  nr02d0 U70 ( .A1(n45), .A2(n27), .ZN(n93) );
  nr02d0 U71 ( .A1(n46), .A2(n27), .ZN(n94) );
  nr02d0 U72 ( .A1(n47), .A2(n27), .ZN(n95) );
  nr02d0 U73 ( .A1(n36), .A2(n28), .ZN(n96) );
  nr02d0 U74 ( .A1(n37), .A2(n28), .ZN(n97) );
  nr02d0 U75 ( .A1(n38), .A2(n28), .ZN(n98) );
  nr02d0 U76 ( .A1(n39), .A2(n28), .ZN(n99) );
  nr02d0 U77 ( .A1(n40), .A2(n28), .ZN(n100) );
  nr02d0 U78 ( .A1(n41), .A2(n28), .ZN(n101) );
  nr02d0 U79 ( .A1(n42), .A2(n28), .ZN(n102) );
  nr02d0 U80 ( .A1(n43), .A2(n28), .ZN(n103) );
  nr02d0 U81 ( .A1(n44), .A2(n28), .ZN(n104) );
  nr02d0 U82 ( .A1(n45), .A2(n28), .ZN(n105) );
  nr02d0 U83 ( .A1(n46), .A2(n28), .ZN(n106) );
  nr02d0 U84 ( .A1(n47), .A2(n28), .ZN(n107) );
  nr02d0 U85 ( .A1(n36), .A2(n29), .ZN(n108) );
  nr02d0 U86 ( .A1(n37), .A2(n29), .ZN(n109) );
  nr02d0 U87 ( .A1(n38), .A2(n29), .ZN(n110) );
  nr02d0 U88 ( .A1(n39), .A2(n29), .ZN(n111) );
  nr02d0 U89 ( .A1(n40), .A2(n29), .ZN(n112) );
  nr02d0 U90 ( .A1(n41), .A2(n29), .ZN(n113) );
  nr02d0 U91 ( .A1(n42), .A2(n29), .ZN(n114) );
  nr02d0 U92 ( .A1(n43), .A2(n29), .ZN(n115) );
  nr02d0 U93 ( .A1(n44), .A2(n29), .ZN(n116) );
  nr02d0 U94 ( .A1(n45), .A2(n29), .ZN(n117) );
  nr02d0 U95 ( .A1(n46), .A2(n29), .ZN(n118) );
  nr02d0 U96 ( .A1(n47), .A2(n29), .ZN(n119) );
  nr02d0 U97 ( .A1(n36), .A2(n30), .ZN(n120) );
  nr02d0 U98 ( .A1(n37), .A2(n30), .ZN(n121) );
  nr02d0 U99 ( .A1(n38), .A2(n30), .ZN(n122) );
  nr02d0 U100 ( .A1(n39), .A2(n30), .ZN(n123) );
  nr02d0 U101 ( .A1(n40), .A2(n30), .ZN(n124) );
  nr02d0 U102 ( .A1(n41), .A2(n30), .ZN(n125) );
  nr02d0 U103 ( .A1(n42), .A2(n30), .ZN(n126) );
  nr02d0 U104 ( .A1(n43), .A2(n30), .ZN(n127) );
  nr02d0 U105 ( .A1(n44), .A2(n30), .ZN(n128) );
  nr02d0 U106 ( .A1(n45), .A2(n30), .ZN(n129) );
  nr02d0 U107 ( .A1(n46), .A2(n30), .ZN(n130) );
  nr02d0 U108 ( .A1(n47), .A2(n30), .ZN(n131) );
  nr02d0 U109 ( .A1(n36), .A2(n31), .ZN(n132) );
  nr02d0 U110 ( .A1(n37), .A2(n31), .ZN(n133) );
  nr02d0 U111 ( .A1(n38), .A2(n31), .ZN(n134) );
  nr02d0 U112 ( .A1(n39), .A2(n31), .ZN(n135) );
  nr02d0 U113 ( .A1(n40), .A2(n31), .ZN(n136) );
  nr02d0 U114 ( .A1(n41), .A2(n31), .ZN(n137) );
  nr02d0 U115 ( .A1(n42), .A2(n31), .ZN(n138) );
  nr02d0 U116 ( .A1(n43), .A2(n31), .ZN(n139) );
  nr02d0 U117 ( .A1(n44), .A2(n31), .ZN(n140) );
  nr02d0 U118 ( .A1(n45), .A2(n31), .ZN(n141) );
  nr02d0 U119 ( .A1(n46), .A2(n31), .ZN(n142) );
  nr02d0 U120 ( .A1(n47), .A2(n31), .ZN(n143) );
  nr02d0 U121 ( .A1(n36), .A2(n32), .ZN(n144) );
  nr02d0 U122 ( .A1(n37), .A2(n32), .ZN(n145) );
  nr02d0 U123 ( .A1(n38), .A2(n32), .ZN(n146) );
  nr02d0 U124 ( .A1(n39), .A2(n32), .ZN(n147) );
  nr02d0 U125 ( .A1(n40), .A2(n32), .ZN(n148) );
  nr02d0 U126 ( .A1(n41), .A2(n32), .ZN(n149) );
  nr02d0 U127 ( .A1(n42), .A2(n32), .ZN(n150) );
  nr02d0 U128 ( .A1(n43), .A2(n32), .ZN(n151) );
  nr02d0 U129 ( .A1(n44), .A2(n32), .ZN(n152) );
  nr02d0 U130 ( .A1(n45), .A2(n32), .ZN(n153) );
  nr02d0 U131 ( .A1(n46), .A2(n32), .ZN(n154) );
  nr02d0 U132 ( .A1(n47), .A2(n32), .ZN(n155) );
  nr02d0 U133 ( .A1(n36), .A2(n33), .ZN(n156) );
  nr02d0 U134 ( .A1(n37), .A2(n33), .ZN(n157) );
  nr02d0 U135 ( .A1(n38), .A2(n33), .ZN(n158) );
  nr02d0 U136 ( .A1(n39), .A2(n33), .ZN(n159) );
  nr02d0 U137 ( .A1(n40), .A2(n33), .ZN(n160) );
  nr02d0 U138 ( .A1(n41), .A2(n33), .ZN(n161) );
  nr02d0 U139 ( .A1(n42), .A2(n33), .ZN(n162) );
  nr02d0 U140 ( .A1(n43), .A2(n33), .ZN(n163) );
  nr02d0 U141 ( .A1(n44), .A2(n33), .ZN(n164) );
  nr02d0 U142 ( .A1(n45), .A2(n33), .ZN(n165) );
  nr02d0 U143 ( .A1(n46), .A2(n33), .ZN(n166) );
  nr02d0 U144 ( .A1(n47), .A2(n33), .ZN(n167) );
  nr02d0 U145 ( .A1(n36), .A2(n34), .ZN(n168) );
  nr02d0 U146 ( .A1(n37), .A2(n34), .ZN(n169) );
  nr02d0 U147 ( .A1(n38), .A2(n34), .ZN(n170) );
  nr02d0 U148 ( .A1(n39), .A2(n34), .ZN(n171) );
  nr02d0 U149 ( .A1(n40), .A2(n34), .ZN(n172) );
  nr02d0 U150 ( .A1(n41), .A2(n34), .ZN(n173) );
  nr02d0 U151 ( .A1(n42), .A2(n34), .ZN(n174) );
  nr02d0 U152 ( .A1(n43), .A2(n34), .ZN(n175) );
  nr02d0 U153 ( .A1(n44), .A2(n34), .ZN(n176) );
  nr02d0 U154 ( .A1(n45), .A2(n34), .ZN(n177) );
  nr02d0 U155 ( .A1(n46), .A2(n34), .ZN(n178) );
  nr02d0 U156 ( .A1(n47), .A2(n34), .ZN(n179) );
  nr02d0 U157 ( .A1(n36), .A2(n35), .ZN(n180) );
  nr02d0 U158 ( .A1(n37), .A2(n35), .ZN(n181) );
  nr02d0 U159 ( .A1(n38), .A2(n35), .ZN(n182) );
  nr02d0 U160 ( .A1(n39), .A2(n35), .ZN(n183) );
  nr02d0 U161 ( .A1(n40), .A2(n35), .ZN(n184) );
  nr02d0 U162 ( .A1(n41), .A2(n35), .ZN(n185) );
  nr02d0 U163 ( .A1(n42), .A2(n35), .ZN(n186) );
  nr02d0 U164 ( .A1(n43), .A2(n35), .ZN(n187) );
  nr02d0 U165 ( .A1(n44), .A2(n35), .ZN(n188) );
  nr02d0 U166 ( .A1(n45), .A2(n35), .ZN(n189) );
  nr02d0 U167 ( .A1(n46), .A2(n35), .ZN(n190) );
  nr02d0 U168 ( .A1(n47), .A2(n35), .ZN(n191) );
  ah01d0 U169 ( .A(n50), .B(n61), .CO(n193), .S(n192) );
  ah01d0 U170 ( .A(n73), .B(n84), .CO(n195), .S(n194) );
  ad01d0 U171 ( .A(n51), .B(n62), .CI(n193), .CO(n197), .S(n196) );
  ah01d0 U172 ( .A(n85), .B(n96), .CO(n199), .S(n198) );
  ad01d0 U173 ( .A(n52), .B(n74), .CI(n63), .CO(n201), .S(n200) );
  ad01d0 U174 ( .A(n195), .B(n198), .CI(n200), .CO(n203), .S(n202) );
  ah01d0 U175 ( .A(n97), .B(n108), .CO(n205), .S(n204) );
  ad01d0 U176 ( .A(n53), .B(n86), .CI(n75), .CO(n207), .S(n206) );
  ad01d0 U177 ( .A(n64), .B(n199), .CI(n204), .CO(n209), .S(n208) );
  ad01d0 U178 ( .A(n201), .B(n206), .CI(n208), .CO(n211), .S(n210) );
  ah01d0 U179 ( .A(n109), .B(n120), .CO(n213), .S(n212) );
  ad01d0 U180 ( .A(n54), .B(n98), .CI(n65), .CO(n215), .S(n214) );
  ad01d0 U181 ( .A(n76), .B(n87), .CI(n205), .CO(n217), .S(n216) );
  ad01d0 U182 ( .A(n212), .B(n207), .CI(n214), .CO(n219), .S(n218) );
  ad01d0 U183 ( .A(n209), .B(n216), .CI(n218), .CO(n221), .S(n220) );
  ah01d0 U184 ( .A(n121), .B(n132), .CO(n223), .S(n222) );
  ad01d0 U185 ( .A(n55), .B(n110), .CI(n66), .CO(n225), .S(n224) );
  ad01d0 U186 ( .A(n77), .B(n99), .CI(n88), .CO(n227), .S(n226) );
  ad01d0 U187 ( .A(n213), .B(n222), .CI(n215), .CO(n229), .S(n228) );
  ad01d0 U188 ( .A(n226), .B(n224), .CI(n217), .CO(n231), .S(n230) );
  ad01d0 U189 ( .A(n228), .B(n219), .CI(n230), .CO(n233), .S(n232) );
  ah01d0 U190 ( .A(n133), .B(n144), .CO(n235), .S(n234) );
  ad01d0 U191 ( .A(n56), .B(n122), .CI(n67), .CO(n237), .S(n236) );
  ad01d0 U192 ( .A(n100), .B(n78), .CI(n111), .CO(n239), .S(n238) );
  ad01d0 U193 ( .A(n89), .B(n223), .CI(n234), .CO(n241), .S(n240) );
  ad01d0 U194 ( .A(n225), .B(n227), .CI(n238), .CO(n243), .S(n242) );
  ad01d0 U195 ( .A(n236), .B(n229), .CI(n240), .CO(n245), .S(n244) );
  ad01d0 U196 ( .A(n231), .B(n242), .CI(n244), .CO(n247), .S(n246) );
  ah01d0 U197 ( .A(n145), .B(n156), .CO(n249), .S(n248) );
  ad01d0 U198 ( .A(n57), .B(n134), .CI(n68), .CO(n251), .S(n250) );
  ad01d0 U199 ( .A(n112), .B(n123), .CI(n101), .CO(n253), .S(n252) );
  ad01d0 U200 ( .A(n79), .B(n90), .CI(n235), .CO(n255), .S(n254) );
  ad01d0 U201 ( .A(n248), .B(n237), .CI(n239), .CO(n257), .S(n256) );
  ad01d0 U202 ( .A(n252), .B(n250), .CI(n241), .CO(n259), .S(n258) );
  ad01d0 U203 ( .A(n254), .B(n243), .CI(n256), .CO(n261), .S(n260) );
  ad01d0 U204 ( .A(n258), .B(n245), .CI(n260), .CO(n263), .S(n262) );
  ah01d0 U205 ( .A(n157), .B(n168), .CO(n265), .S(n264) );
  ad01d0 U206 ( .A(n58), .B(n146), .CI(n135), .CO(n267), .S(n266) );
  ad01d0 U207 ( .A(n102), .B(n69), .CI(n124), .CO(n269), .S(n268) );
  ad01d0 U208 ( .A(n80), .B(n113), .CI(n91), .CO(n271), .S(n270) );
  ad01d0 U209 ( .A(n249), .B(n264), .CI(n251), .CO(n273), .S(n272) );
  ad01d0 U210 ( .A(n253), .B(n270), .CI(n268), .CO(n275), .S(n274) );
  ad01d0 U211 ( .A(n266), .B(n255), .CI(n257), .CO(n277), .S(n276) );
  ad01d0 U212 ( .A(n272), .B(n259), .CI(n274), .CO(n279), .S(n278) );
  ad01d0 U213 ( .A(n276), .B(n261), .CI(n278), .CO(n281), .S(n280) );
  ah01d0 U214 ( .A(n169), .B(n180), .CO(n283), .S(n282) );
  ad01d0 U215 ( .A(n59), .B(n158), .CI(n70), .CO(n285), .S(n284) );
  ad01d0 U216 ( .A(n125), .B(n147), .CI(n136), .CO(n287), .S(n286) );
  ad01d0 U217 ( .A(n81), .B(n114), .CI(n103), .CO(n289), .S(n288) );
  ad01d0 U218 ( .A(n92), .B(n265), .CI(n282), .CO(n291), .S(n290) );
  ad01d0 U219 ( .A(n267), .B(n271), .CI(n269), .CO(n293), .S(n292) );
  ad01d0 U220 ( .A(n288), .B(n284), .CI(n286), .CO(n295), .S(n294) );
  ad01d0 U221 ( .A(n273), .B(n290), .CI(n275), .CO(n297), .S(n296) );
  ad01d0 U222 ( .A(n292), .B(n294), .CI(n277), .CO(n299), .S(n298) );
  ad01d0 U223 ( .A(n296), .B(n279), .CI(n298), .CO(n301), .S(n300) );
  ah01d0 U224 ( .A(n170), .B(n181), .CO(n303), .S(n302) );
  ad01d0 U225 ( .A(n126), .B(n71), .CI(n82), .CO(n305), .S(n304) );
  ad01d0 U226 ( .A(n137), .B(n159), .CI(n148), .CO(n307), .S(n306) );
  ad01d0 U227 ( .A(n93), .B(n115), .CI(n104), .CO(n309), .S(n308) );
  ad01d0 U228 ( .A(n283), .B(n302), .CI(n285), .CO(n311), .S(n310) );
  ad01d0 U229 ( .A(n287), .B(n289), .CI(n308), .CO(n313), .S(n312) );
  ad01d0 U230 ( .A(n306), .B(n304), .CI(n291), .CO(n315), .S(n314) );
  ad01d0 U231 ( .A(n293), .B(n310), .CI(n295), .CO(n317), .S(n316) );
  ad01d0 U232 ( .A(n312), .B(n314), .CI(n297), .CO(n319), .S(n318) );
  ad01d0 U233 ( .A(n316), .B(n299), .CI(n318), .CO(n321), .S(n320) );
  ad01d0 U234 ( .A(n83), .B(n182), .CI(n171), .CO(n323), .S(n322) );
  ad01d0 U235 ( .A(n94), .B(n160), .CI(n149), .CO(n325), .S(n324) );
  ad01d0 U236 ( .A(n105), .B(n138), .CI(n127), .CO(n327), .S(n326) );
  ad01d0 U237 ( .A(n116), .B(n303), .CI(n305), .CO(n329), .S(n328) );
  ad01d0 U238 ( .A(n307), .B(n309), .CI(n326), .CO(n331), .S(n330) );
  ad01d0 U239 ( .A(n324), .B(n322), .CI(n311), .CO(n333), .S(n332) );
  ad01d0 U240 ( .A(n328), .B(n313), .CI(n315), .CO(n335), .S(n334) );
  ad01d0 U241 ( .A(n330), .B(n332), .CI(n317), .CO(n337), .S(n336) );
  ad01d0 U242 ( .A(n334), .B(n319), .CI(n336), .CO(n339), .S(n338) );
  ad01d0 U243 ( .A(n95), .B(n183), .CI(n172), .CO(n341), .S(n340) );
  ad01d0 U244 ( .A(n106), .B(n161), .CI(n117), .CO(n343), .S(n342) );
  ad01d0 U245 ( .A(n128), .B(n150), .CI(n139), .CO(n345), .S(n344) );
  ad01d0 U246 ( .A(n323), .B(n327), .CI(n325), .CO(n347), .S(n346) );
  ad01d0 U247 ( .A(n344), .B(n340), .CI(n342), .CO(n349), .S(n348) );
  ad01d0 U248 ( .A(n329), .B(n331), .CI(n346), .CO(n351), .S(n350) );
  ad01d0 U249 ( .A(n333), .B(n348), .CI(n335), .CO(n353), .S(n352) );
  ad01d0 U250 ( .A(n350), .B(n337), .CI(n352), .CO(n355), .S(n354) );
  ad01d0 U251 ( .A(n107), .B(n184), .CI(n173), .CO(n357), .S(n356) );
  ad01d0 U252 ( .A(n118), .B(n162), .CI(n151), .CO(n359), .S(n358) );
  ad01d0 U253 ( .A(n129), .B(n140), .CI(n341), .CO(n361), .S(n360) );
  ad01d0 U254 ( .A(n343), .B(n345), .CI(n358), .CO(n363), .S(n362) );
  ad01d0 U255 ( .A(n356), .B(n347), .CI(n360), .CO(n365), .S(n364) );
  ad01d0 U256 ( .A(n349), .B(n362), .CI(n351), .CO(n367), .S(n366) );
  ad01d0 U257 ( .A(n364), .B(n353), .CI(n366), .CO(n369), .S(n368) );
  ad01d0 U258 ( .A(n119), .B(n185), .CI(n174), .CO(n371), .S(n370) );
  ad01d0 U259 ( .A(n163), .B(n130), .CI(n141), .CO(n373), .S(n372) );
  ad01d0 U260 ( .A(n152), .B(n357), .CI(n359), .CO(n375), .S(n374) );
  ad01d0 U261 ( .A(n372), .B(n370), .CI(n361), .CO(n377), .S(n376) );
  ad01d0 U262 ( .A(n363), .B(n374), .CI(n376), .CO(n379), .S(n378) );
  ad01d0 U263 ( .A(n365), .B(n367), .CI(n378), .CO(n381), .S(n380) );
  ad01d0 U264 ( .A(n131), .B(n186), .CI(n175), .CO(n383), .S(n382) );
  ad01d0 U265 ( .A(n164), .B(n153), .CI(n142), .CO(n385), .S(n384) );
  ad01d0 U266 ( .A(n371), .B(n373), .CI(n384), .CO(n387), .S(n386) );
  ad01d0 U267 ( .A(n382), .B(n375), .CI(n386), .CO(n389), .S(n388) );
  ad01d0 U268 ( .A(n377), .B(n388), .CI(n379), .CO(n391), .S(n390) );
  ad01d0 U269 ( .A(n143), .B(n187), .CI(n176), .CO(n393), .S(n392) );
  ad01d0 U270 ( .A(n154), .B(n165), .CI(n383), .CO(n395), .S(n394) );
  ad01d0 U271 ( .A(n385), .B(n392), .CI(n394), .CO(n397), .S(n396) );
  ad01d0 U272 ( .A(n387), .B(n396), .CI(n389), .CO(n399), .S(n398) );
  ad01d0 U273 ( .A(n155), .B(n188), .CI(n177), .CO(n401), .S(n400) );
  ad01d0 U274 ( .A(n166), .B(n393), .CI(n400), .CO(n403), .S(n402) );
  ad01d0 U275 ( .A(n395), .B(n402), .CI(n397), .CO(n405), .S(n404) );
  ad01d0 U276 ( .A(n167), .B(n189), .CI(n178), .CO(n407), .S(n406) );
  ad01d0 U277 ( .A(n401), .B(n406), .CI(n403), .CO(n409), .S(n408) );
  ad01d0 U278 ( .A(n179), .B(n190), .CI(n407), .CO(n411), .S(n410) );
  ah01d0 U279 ( .A(n60), .B(n49), .CO(n412), .S(product[1]) );
  ad01d0 U280 ( .A(n72), .B(n412), .CI(n192), .CO(n413), .S(product[2]) );
  ad01d0 U281 ( .A(n194), .B(n413), .CI(n196), .CO(n414), .S(product[3]) );
  ad01d0 U282 ( .A(n197), .B(n202), .CI(n414), .CO(n415), .S(product[4]) );
  ad01d0 U283 ( .A(n203), .B(n210), .CI(n415), .CO(n416), .S(product[5]) );
  ad01d0 U284 ( .A(n211), .B(n220), .CI(n416), .CO(n417), .S(product[6]) );
  ad01d0 U285 ( .A(n221), .B(n232), .CI(n417), .CO(n418), .S(product[7]) );
  ad01d0 U286 ( .A(n233), .B(n246), .CI(n418), .CO(n419), .S(product[8]) );
  ad01d0 U287 ( .A(n247), .B(n262), .CI(n419), .CO(n420), .S(product[9]) );
  ad01d0 U288 ( .A(n263), .B(n280), .CI(n420), .CO(n421), .S(product[10]) );
  ad01d0 U289 ( .A(n281), .B(n300), .CI(n421), .CO(n422), .S(product[11]) );
  ad01d0 U290 ( .A(n301), .B(n320), .CI(n422), .CO(n423), .S(product[12]) );
  ad01d0 U291 ( .A(n321), .B(n338), .CI(n423), .CO(n424), .S(product[13]) );
  ad01d0 U292 ( .A(n339), .B(n354), .CI(n424), .CO(n425), .S(product[14]) );
  ad01d0 U295 ( .A(n390), .B(n381), .CI(n427), .CO(n428), .S(product[17]) );
  ad01d0 U296 ( .A(n398), .B(n391), .CI(n428), .CO(n429), .S(product[18]) );
  ad01d0 U297 ( .A(n404), .B(n399), .CI(n429), .CO(n430), .S(product[19]) );
  ad01d0 U298 ( .A(n408), .B(n405), .CI(n430), .CO(n431), .S(product[20]) );
  ad01d0 U299 ( .A(n410), .B(n409), .CI(n431), .CO(n432), .S(product[21]) );
  ad01d0 U300 ( .A(n191), .B(n411), .CI(n432), .CO(product[23]), .S(
        product[22]) );
  ad01d0 U304 ( .A(n355), .B(n368), .CI(n425), .CO(n426), .S(product[15]) );
  ad01d0 U305 ( .A(n369), .B(n380), .CI(n426), .CO(n427), .S(product[16]) );
  inv0d1 U306 ( .I(b[3]), .ZN(n39) );
  inv0d1 U307 ( .I(b[4]), .ZN(n40) );
  inv0d1 U308 ( .I(b[5]), .ZN(n41) );
  inv0d1 U309 ( .I(b[6]), .ZN(n42) );
  inv0d1 U310 ( .I(b[0]), .ZN(n36) );
  inv0d1 U311 ( .I(b[1]), .ZN(n37) );
  inv0d1 U312 ( .I(a[0]), .ZN(n24) );
  inv0d1 U313 ( .I(a[3]), .ZN(n27) );
  inv0d1 U314 ( .I(a[5]), .ZN(n29) );
  inv0d1 U315 ( .I(a[4]), .ZN(n28) );
  inv0d1 U316 ( .I(a[1]), .ZN(n25) );
  inv0d1 U317 ( .I(a[2]), .ZN(n26) );
  inv0d1 U318 ( .I(b[2]), .ZN(n38) );
  inv0d1 U319 ( .I(b[7]), .ZN(n43) );
  inv0d1 U320 ( .I(a[6]), .ZN(n30) );
  inv0d1 U321 ( .I(a[7]), .ZN(n31) );
  inv0d1 U322 ( .I(a[8]), .ZN(n32) );
  inv0d1 U323 ( .I(a[9]), .ZN(n33) );
  inv0d1 U324 ( .I(a[10]), .ZN(n34) );
  inv0d1 U325 ( .I(b[8]), .ZN(n44) );
  inv0d1 U326 ( .I(b[10]), .ZN(n46) );
  inv0d1 U327 ( .I(b[11]), .ZN(n47) );
  inv0d1 U328 ( .I(b[9]), .ZN(n45) );
  inv0d1 U329 ( .I(a[11]), .ZN(n35) );
endmodule


module BLENDER_DW_mult_uns_4 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432;

  nr02d0 U25 ( .A1(n36), .A2(n24), .ZN(product[0]) );
  nr02d0 U26 ( .A1(n37), .A2(n24), .ZN(n49) );
  nr02d0 U27 ( .A1(n38), .A2(n24), .ZN(n50) );
  nr02d0 U28 ( .A1(n39), .A2(n24), .ZN(n51) );
  nr02d0 U29 ( .A1(n40), .A2(n24), .ZN(n52) );
  nr02d0 U30 ( .A1(n41), .A2(n24), .ZN(n53) );
  nr02d0 U31 ( .A1(n42), .A2(n24), .ZN(n54) );
  nr02d0 U32 ( .A1(n43), .A2(n24), .ZN(n55) );
  nr02d0 U33 ( .A1(n44), .A2(n24), .ZN(n56) );
  nr02d0 U34 ( .A1(n45), .A2(n24), .ZN(n57) );
  nr02d0 U35 ( .A1(n46), .A2(n24), .ZN(n58) );
  nr02d0 U36 ( .A1(n47), .A2(n24), .ZN(n59) );
  nr02d0 U37 ( .A1(n36), .A2(n25), .ZN(n60) );
  nr02d0 U38 ( .A1(n37), .A2(n25), .ZN(n61) );
  nr02d0 U39 ( .A1(n38), .A2(n25), .ZN(n62) );
  nr02d0 U40 ( .A1(n39), .A2(n25), .ZN(n63) );
  nr02d0 U41 ( .A1(n40), .A2(n25), .ZN(n64) );
  nr02d0 U42 ( .A1(n41), .A2(n25), .ZN(n65) );
  nr02d0 U43 ( .A1(n42), .A2(n25), .ZN(n66) );
  nr02d0 U44 ( .A1(n43), .A2(n25), .ZN(n67) );
  nr02d0 U45 ( .A1(n44), .A2(n25), .ZN(n68) );
  nr02d0 U46 ( .A1(n45), .A2(n25), .ZN(n69) );
  nr02d0 U47 ( .A1(n46), .A2(n25), .ZN(n70) );
  nr02d0 U48 ( .A1(n47), .A2(n25), .ZN(n71) );
  nr02d0 U49 ( .A1(n36), .A2(n26), .ZN(n72) );
  nr02d0 U50 ( .A1(n37), .A2(n26), .ZN(n73) );
  nr02d0 U51 ( .A1(n38), .A2(n26), .ZN(n74) );
  nr02d0 U52 ( .A1(n39), .A2(n26), .ZN(n75) );
  nr02d0 U53 ( .A1(n40), .A2(n26), .ZN(n76) );
  nr02d0 U54 ( .A1(n41), .A2(n26), .ZN(n77) );
  nr02d0 U55 ( .A1(n42), .A2(n26), .ZN(n78) );
  nr02d0 U56 ( .A1(n43), .A2(n26), .ZN(n79) );
  nr02d0 U57 ( .A1(n44), .A2(n26), .ZN(n80) );
  nr02d0 U58 ( .A1(n45), .A2(n26), .ZN(n81) );
  nr02d0 U59 ( .A1(n46), .A2(n26), .ZN(n82) );
  nr02d0 U60 ( .A1(n47), .A2(n26), .ZN(n83) );
  nr02d0 U61 ( .A1(n36), .A2(n27), .ZN(n84) );
  nr02d0 U62 ( .A1(n37), .A2(n27), .ZN(n85) );
  nr02d0 U63 ( .A1(n38), .A2(n27), .ZN(n86) );
  nr02d0 U64 ( .A1(n39), .A2(n27), .ZN(n87) );
  nr02d0 U65 ( .A1(n40), .A2(n27), .ZN(n88) );
  nr02d0 U66 ( .A1(n41), .A2(n27), .ZN(n89) );
  nr02d0 U67 ( .A1(n42), .A2(n27), .ZN(n90) );
  nr02d0 U68 ( .A1(n43), .A2(n27), .ZN(n91) );
  nr02d0 U69 ( .A1(n44), .A2(n27), .ZN(n92) );
  nr02d0 U70 ( .A1(n45), .A2(n27), .ZN(n93) );
  nr02d0 U71 ( .A1(n46), .A2(n27), .ZN(n94) );
  nr02d0 U72 ( .A1(n47), .A2(n27), .ZN(n95) );
  nr02d0 U73 ( .A1(n36), .A2(n28), .ZN(n96) );
  nr02d0 U74 ( .A1(n37), .A2(n28), .ZN(n97) );
  nr02d0 U75 ( .A1(n38), .A2(n28), .ZN(n98) );
  nr02d0 U76 ( .A1(n39), .A2(n28), .ZN(n99) );
  nr02d0 U77 ( .A1(n40), .A2(n28), .ZN(n100) );
  nr02d0 U78 ( .A1(n41), .A2(n28), .ZN(n101) );
  nr02d0 U79 ( .A1(n42), .A2(n28), .ZN(n102) );
  nr02d0 U80 ( .A1(n43), .A2(n28), .ZN(n103) );
  nr02d0 U81 ( .A1(n44), .A2(n28), .ZN(n104) );
  nr02d0 U82 ( .A1(n45), .A2(n28), .ZN(n105) );
  nr02d0 U83 ( .A1(n46), .A2(n28), .ZN(n106) );
  nr02d0 U84 ( .A1(n47), .A2(n28), .ZN(n107) );
  nr02d0 U85 ( .A1(n36), .A2(n29), .ZN(n108) );
  nr02d0 U86 ( .A1(n37), .A2(n29), .ZN(n109) );
  nr02d0 U87 ( .A1(n38), .A2(n29), .ZN(n110) );
  nr02d0 U88 ( .A1(n39), .A2(n29), .ZN(n111) );
  nr02d0 U89 ( .A1(n40), .A2(n29), .ZN(n112) );
  nr02d0 U90 ( .A1(n41), .A2(n29), .ZN(n113) );
  nr02d0 U91 ( .A1(n42), .A2(n29), .ZN(n114) );
  nr02d0 U92 ( .A1(n43), .A2(n29), .ZN(n115) );
  nr02d0 U93 ( .A1(n44), .A2(n29), .ZN(n116) );
  nr02d0 U94 ( .A1(n45), .A2(n29), .ZN(n117) );
  nr02d0 U95 ( .A1(n46), .A2(n29), .ZN(n118) );
  nr02d0 U96 ( .A1(n47), .A2(n29), .ZN(n119) );
  nr02d0 U97 ( .A1(n36), .A2(n30), .ZN(n120) );
  nr02d0 U98 ( .A1(n37), .A2(n30), .ZN(n121) );
  nr02d0 U99 ( .A1(n38), .A2(n30), .ZN(n122) );
  nr02d0 U100 ( .A1(n39), .A2(n30), .ZN(n123) );
  nr02d0 U101 ( .A1(n40), .A2(n30), .ZN(n124) );
  nr02d0 U102 ( .A1(n41), .A2(n30), .ZN(n125) );
  nr02d0 U103 ( .A1(n42), .A2(n30), .ZN(n126) );
  nr02d0 U104 ( .A1(n43), .A2(n30), .ZN(n127) );
  nr02d0 U105 ( .A1(n44), .A2(n30), .ZN(n128) );
  nr02d0 U106 ( .A1(n45), .A2(n30), .ZN(n129) );
  nr02d0 U107 ( .A1(n46), .A2(n30), .ZN(n130) );
  nr02d0 U108 ( .A1(n47), .A2(n30), .ZN(n131) );
  nr02d0 U109 ( .A1(n36), .A2(n31), .ZN(n132) );
  nr02d0 U110 ( .A1(n37), .A2(n31), .ZN(n133) );
  nr02d0 U111 ( .A1(n38), .A2(n31), .ZN(n134) );
  nr02d0 U112 ( .A1(n39), .A2(n31), .ZN(n135) );
  nr02d0 U113 ( .A1(n40), .A2(n31), .ZN(n136) );
  nr02d0 U114 ( .A1(n41), .A2(n31), .ZN(n137) );
  nr02d0 U115 ( .A1(n42), .A2(n31), .ZN(n138) );
  nr02d0 U116 ( .A1(n43), .A2(n31), .ZN(n139) );
  nr02d0 U117 ( .A1(n44), .A2(n31), .ZN(n140) );
  nr02d0 U118 ( .A1(n45), .A2(n31), .ZN(n141) );
  nr02d0 U119 ( .A1(n46), .A2(n31), .ZN(n142) );
  nr02d0 U120 ( .A1(n47), .A2(n31), .ZN(n143) );
  nr02d0 U121 ( .A1(n36), .A2(n32), .ZN(n144) );
  nr02d0 U122 ( .A1(n37), .A2(n32), .ZN(n145) );
  nr02d0 U123 ( .A1(n38), .A2(n32), .ZN(n146) );
  nr02d0 U124 ( .A1(n39), .A2(n32), .ZN(n147) );
  nr02d0 U125 ( .A1(n40), .A2(n32), .ZN(n148) );
  nr02d0 U126 ( .A1(n41), .A2(n32), .ZN(n149) );
  nr02d0 U127 ( .A1(n42), .A2(n32), .ZN(n150) );
  nr02d0 U128 ( .A1(n43), .A2(n32), .ZN(n151) );
  nr02d0 U129 ( .A1(n44), .A2(n32), .ZN(n152) );
  nr02d0 U130 ( .A1(n45), .A2(n32), .ZN(n153) );
  nr02d0 U131 ( .A1(n46), .A2(n32), .ZN(n154) );
  nr02d0 U132 ( .A1(n47), .A2(n32), .ZN(n155) );
  nr02d0 U133 ( .A1(n36), .A2(n33), .ZN(n156) );
  nr02d0 U134 ( .A1(n37), .A2(n33), .ZN(n157) );
  nr02d0 U135 ( .A1(n38), .A2(n33), .ZN(n158) );
  nr02d0 U136 ( .A1(n39), .A2(n33), .ZN(n159) );
  nr02d0 U137 ( .A1(n40), .A2(n33), .ZN(n160) );
  nr02d0 U138 ( .A1(n41), .A2(n33), .ZN(n161) );
  nr02d0 U139 ( .A1(n42), .A2(n33), .ZN(n162) );
  nr02d0 U140 ( .A1(n43), .A2(n33), .ZN(n163) );
  nr02d0 U141 ( .A1(n44), .A2(n33), .ZN(n164) );
  nr02d0 U142 ( .A1(n45), .A2(n33), .ZN(n165) );
  nr02d0 U143 ( .A1(n46), .A2(n33), .ZN(n166) );
  nr02d0 U144 ( .A1(n47), .A2(n33), .ZN(n167) );
  nr02d0 U145 ( .A1(n36), .A2(n34), .ZN(n168) );
  nr02d0 U146 ( .A1(n37), .A2(n34), .ZN(n169) );
  nr02d0 U147 ( .A1(n38), .A2(n34), .ZN(n170) );
  nr02d0 U148 ( .A1(n39), .A2(n34), .ZN(n171) );
  nr02d0 U149 ( .A1(n40), .A2(n34), .ZN(n172) );
  nr02d0 U150 ( .A1(n41), .A2(n34), .ZN(n173) );
  nr02d0 U151 ( .A1(n42), .A2(n34), .ZN(n174) );
  nr02d0 U152 ( .A1(n43), .A2(n34), .ZN(n175) );
  nr02d0 U153 ( .A1(n44), .A2(n34), .ZN(n176) );
  nr02d0 U154 ( .A1(n45), .A2(n34), .ZN(n177) );
  nr02d0 U155 ( .A1(n46), .A2(n34), .ZN(n178) );
  nr02d0 U156 ( .A1(n47), .A2(n34), .ZN(n179) );
  nr02d0 U157 ( .A1(n36), .A2(n35), .ZN(n180) );
  nr02d0 U158 ( .A1(n37), .A2(n35), .ZN(n181) );
  nr02d0 U159 ( .A1(n38), .A2(n35), .ZN(n182) );
  nr02d0 U160 ( .A1(n39), .A2(n35), .ZN(n183) );
  nr02d0 U161 ( .A1(n40), .A2(n35), .ZN(n184) );
  nr02d0 U162 ( .A1(n41), .A2(n35), .ZN(n185) );
  nr02d0 U163 ( .A1(n42), .A2(n35), .ZN(n186) );
  nr02d0 U164 ( .A1(n43), .A2(n35), .ZN(n187) );
  nr02d0 U165 ( .A1(n44), .A2(n35), .ZN(n188) );
  nr02d0 U166 ( .A1(n45), .A2(n35), .ZN(n189) );
  nr02d0 U167 ( .A1(n46), .A2(n35), .ZN(n190) );
  nr02d0 U168 ( .A1(n47), .A2(n35), .ZN(n191) );
  ah01d0 U170 ( .A(n73), .B(n84), .CO(n195), .S(n194) );
  ad01d0 U171 ( .A(n51), .B(n62), .CI(n193), .CO(n197), .S(n196) );
  ah01d0 U172 ( .A(n85), .B(n96), .CO(n199), .S(n198) );
  ad01d0 U173 ( .A(n52), .B(n74), .CI(n63), .CO(n201), .S(n200) );
  ad01d0 U174 ( .A(n195), .B(n198), .CI(n200), .CO(n203), .S(n202) );
  ah01d0 U175 ( .A(n97), .B(n108), .CO(n205), .S(n204) );
  ad01d0 U176 ( .A(n53), .B(n86), .CI(n75), .CO(n207), .S(n206) );
  ad01d0 U177 ( .A(n64), .B(n199), .CI(n204), .CO(n209), .S(n208) );
  ad01d0 U178 ( .A(n201), .B(n206), .CI(n208), .CO(n211), .S(n210) );
  ah01d0 U179 ( .A(n109), .B(n120), .CO(n213), .S(n212) );
  ad01d0 U180 ( .A(n54), .B(n98), .CI(n65), .CO(n215), .S(n214) );
  ad01d0 U181 ( .A(n76), .B(n87), .CI(n205), .CO(n217), .S(n216) );
  ad01d0 U182 ( .A(n212), .B(n207), .CI(n214), .CO(n219), .S(n218) );
  ad01d0 U183 ( .A(n209), .B(n216), .CI(n218), .CO(n221), .S(n220) );
  ah01d0 U184 ( .A(n121), .B(n132), .CO(n223), .S(n222) );
  ad01d0 U185 ( .A(n55), .B(n110), .CI(n66), .CO(n225), .S(n224) );
  ad01d0 U186 ( .A(n77), .B(n99), .CI(n88), .CO(n227), .S(n226) );
  ad01d0 U187 ( .A(n213), .B(n222), .CI(n215), .CO(n229), .S(n228) );
  ad01d0 U188 ( .A(n226), .B(n224), .CI(n217), .CO(n231), .S(n230) );
  ad01d0 U189 ( .A(n228), .B(n219), .CI(n230), .CO(n233), .S(n232) );
  ah01d0 U190 ( .A(n133), .B(n144), .CO(n235), .S(n234) );
  ad01d0 U191 ( .A(n56), .B(n122), .CI(n67), .CO(n237), .S(n236) );
  ad01d0 U192 ( .A(n100), .B(n78), .CI(n111), .CO(n239), .S(n238) );
  ad01d0 U193 ( .A(n89), .B(n223), .CI(n234), .CO(n241), .S(n240) );
  ad01d0 U194 ( .A(n225), .B(n227), .CI(n238), .CO(n243), .S(n242) );
  ad01d0 U195 ( .A(n236), .B(n229), .CI(n240), .CO(n245), .S(n244) );
  ad01d0 U196 ( .A(n231), .B(n242), .CI(n244), .CO(n247), .S(n246) );
  ah01d0 U197 ( .A(n145), .B(n156), .CO(n249), .S(n248) );
  ad01d0 U198 ( .A(n57), .B(n134), .CI(n68), .CO(n251), .S(n250) );
  ad01d0 U199 ( .A(n112), .B(n123), .CI(n101), .CO(n253), .S(n252) );
  ad01d0 U200 ( .A(n79), .B(n90), .CI(n235), .CO(n255), .S(n254) );
  ad01d0 U201 ( .A(n248), .B(n237), .CI(n239), .CO(n257), .S(n256) );
  ad01d0 U202 ( .A(n252), .B(n250), .CI(n241), .CO(n259), .S(n258) );
  ad01d0 U203 ( .A(n254), .B(n243), .CI(n256), .CO(n261), .S(n260) );
  ad01d0 U204 ( .A(n258), .B(n245), .CI(n260), .CO(n263), .S(n262) );
  ah01d0 U205 ( .A(n157), .B(n168), .CO(n265), .S(n264) );
  ad01d0 U206 ( .A(n58), .B(n146), .CI(n135), .CO(n267), .S(n266) );
  ad01d0 U207 ( .A(n102), .B(n69), .CI(n124), .CO(n269), .S(n268) );
  ad01d0 U208 ( .A(n80), .B(n113), .CI(n91), .CO(n271), .S(n270) );
  ad01d0 U209 ( .A(n249), .B(n264), .CI(n251), .CO(n273), .S(n272) );
  ad01d0 U210 ( .A(n253), .B(n270), .CI(n268), .CO(n275), .S(n274) );
  ad01d0 U211 ( .A(n266), .B(n255), .CI(n257), .CO(n277), .S(n276) );
  ad01d0 U212 ( .A(n272), .B(n259), .CI(n274), .CO(n279), .S(n278) );
  ad01d0 U213 ( .A(n276), .B(n261), .CI(n278), .CO(n281), .S(n280) );
  ah01d0 U214 ( .A(n169), .B(n180), .CO(n283), .S(n282) );
  ad01d0 U215 ( .A(n59), .B(n158), .CI(n70), .CO(n285), .S(n284) );
  ad01d0 U216 ( .A(n125), .B(n147), .CI(n136), .CO(n287), .S(n286) );
  ad01d0 U217 ( .A(n81), .B(n114), .CI(n103), .CO(n289), .S(n288) );
  ad01d0 U218 ( .A(n92), .B(n265), .CI(n282), .CO(n291), .S(n290) );
  ad01d0 U219 ( .A(n267), .B(n271), .CI(n269), .CO(n293), .S(n292) );
  ad01d0 U220 ( .A(n288), .B(n284), .CI(n286), .CO(n295), .S(n294) );
  ad01d0 U221 ( .A(n273), .B(n290), .CI(n275), .CO(n297), .S(n296) );
  ad01d0 U222 ( .A(n292), .B(n294), .CI(n277), .CO(n299), .S(n298) );
  ad01d0 U223 ( .A(n296), .B(n279), .CI(n298), .CO(n301), .S(n300) );
  ah01d0 U224 ( .A(n170), .B(n181), .CO(n303), .S(n302) );
  ad01d0 U225 ( .A(n126), .B(n71), .CI(n82), .CO(n305), .S(n304) );
  ad01d0 U226 ( .A(n137), .B(n159), .CI(n148), .CO(n307), .S(n306) );
  ad01d0 U227 ( .A(n93), .B(n115), .CI(n104), .CO(n309), .S(n308) );
  ad01d0 U228 ( .A(n283), .B(n302), .CI(n285), .CO(n311), .S(n310) );
  ad01d0 U229 ( .A(n287), .B(n289), .CI(n308), .CO(n313), .S(n312) );
  ad01d0 U230 ( .A(n306), .B(n304), .CI(n291), .CO(n315), .S(n314) );
  ad01d0 U231 ( .A(n293), .B(n310), .CI(n295), .CO(n317), .S(n316) );
  ad01d0 U232 ( .A(n312), .B(n314), .CI(n297), .CO(n319), .S(n318) );
  ad01d0 U233 ( .A(n316), .B(n299), .CI(n318), .CO(n321), .S(n320) );
  ad01d0 U234 ( .A(n83), .B(n182), .CI(n171), .CO(n323), .S(n322) );
  ad01d0 U235 ( .A(n94), .B(n160), .CI(n149), .CO(n325), .S(n324) );
  ad01d0 U236 ( .A(n105), .B(n138), .CI(n127), .CO(n327), .S(n326) );
  ad01d0 U237 ( .A(n116), .B(n303), .CI(n305), .CO(n329), .S(n328) );
  ad01d0 U238 ( .A(n307), .B(n309), .CI(n326), .CO(n331), .S(n330) );
  ad01d0 U239 ( .A(n324), .B(n322), .CI(n311), .CO(n333), .S(n332) );
  ad01d0 U240 ( .A(n328), .B(n313), .CI(n315), .CO(n335), .S(n334) );
  ad01d0 U241 ( .A(n330), .B(n332), .CI(n317), .CO(n337), .S(n336) );
  ad01d0 U242 ( .A(n334), .B(n319), .CI(n336), .CO(n339), .S(n338) );
  ad01d0 U243 ( .A(n95), .B(n183), .CI(n172), .CO(n341), .S(n340) );
  ad01d0 U244 ( .A(n106), .B(n161), .CI(n117), .CO(n343), .S(n342) );
  ad01d0 U245 ( .A(n128), .B(n150), .CI(n139), .CO(n345), .S(n344) );
  ad01d0 U246 ( .A(n323), .B(n327), .CI(n325), .CO(n347), .S(n346) );
  ad01d0 U247 ( .A(n344), .B(n340), .CI(n342), .CO(n349), .S(n348) );
  ad01d0 U248 ( .A(n329), .B(n331), .CI(n346), .CO(n351), .S(n350) );
  ad01d0 U249 ( .A(n333), .B(n348), .CI(n335), .CO(n353), .S(n352) );
  ad01d0 U250 ( .A(n350), .B(n337), .CI(n352), .CO(n355), .S(n354) );
  ad01d0 U251 ( .A(n107), .B(n184), .CI(n173), .CO(n357), .S(n356) );
  ad01d0 U252 ( .A(n118), .B(n162), .CI(n151), .CO(n359), .S(n358) );
  ad01d0 U253 ( .A(n129), .B(n140), .CI(n341), .CO(n361), .S(n360) );
  ad01d0 U254 ( .A(n343), .B(n345), .CI(n358), .CO(n363), .S(n362) );
  ad01d0 U255 ( .A(n356), .B(n347), .CI(n360), .CO(n365), .S(n364) );
  ad01d0 U256 ( .A(n349), .B(n362), .CI(n351), .CO(n367), .S(n366) );
  ad01d0 U257 ( .A(n364), .B(n353), .CI(n366), .CO(n369), .S(n368) );
  ad01d0 U258 ( .A(n119), .B(n185), .CI(n174), .CO(n371), .S(n370) );
  ad01d0 U259 ( .A(n163), .B(n130), .CI(n141), .CO(n373), .S(n372) );
  ad01d0 U260 ( .A(n152), .B(n357), .CI(n359), .CO(n375), .S(n374) );
  ad01d0 U261 ( .A(n372), .B(n370), .CI(n361), .CO(n377), .S(n376) );
  ad01d0 U262 ( .A(n363), .B(n374), .CI(n376), .CO(n379), .S(n378) );
  ad01d0 U263 ( .A(n365), .B(n367), .CI(n378), .CO(n381), .S(n380) );
  ad01d0 U264 ( .A(n131), .B(n186), .CI(n175), .CO(n383), .S(n382) );
  ad01d0 U265 ( .A(n164), .B(n153), .CI(n142), .CO(n385), .S(n384) );
  ad01d0 U266 ( .A(n371), .B(n373), .CI(n384), .CO(n387), .S(n386) );
  ad01d0 U267 ( .A(n382), .B(n375), .CI(n386), .CO(n389), .S(n388) );
  ad01d0 U268 ( .A(n377), .B(n388), .CI(n379), .CO(n391), .S(n390) );
  ad01d0 U269 ( .A(n143), .B(n187), .CI(n176), .CO(n393), .S(n392) );
  ad01d0 U270 ( .A(n154), .B(n165), .CI(n383), .CO(n395), .S(n394) );
  ad01d0 U271 ( .A(n385), .B(n392), .CI(n394), .CO(n397), .S(n396) );
  ad01d0 U272 ( .A(n387), .B(n396), .CI(n389), .CO(n399), .S(n398) );
  ad01d0 U273 ( .A(n155), .B(n188), .CI(n177), .CO(n401), .S(n400) );
  ad01d0 U274 ( .A(n166), .B(n393), .CI(n400), .CO(n403), .S(n402) );
  ad01d0 U275 ( .A(n395), .B(n402), .CI(n397), .CO(n405), .S(n404) );
  ad01d0 U276 ( .A(n167), .B(n189), .CI(n178), .CO(n407), .S(n406) );
  ad01d0 U277 ( .A(n401), .B(n406), .CI(n403), .CO(n409), .S(n408) );
  ad01d0 U278 ( .A(n179), .B(n190), .CI(n407), .CO(n411), .S(n410) );
  ah01d0 U279 ( .A(n60), .B(n49), .CO(n412), .S(product[1]) );
  ad01d0 U281 ( .A(n194), .B(n413), .CI(n196), .CO(n414), .S(product[3]) );
  ad01d0 U282 ( .A(n197), .B(n202), .CI(n414), .CO(n415), .S(product[4]) );
  ad01d0 U283 ( .A(n203), .B(n210), .CI(n415), .CO(n416), .S(product[5]) );
  ad01d0 U284 ( .A(n211), .B(n220), .CI(n416), .CO(n417), .S(product[6]) );
  ad01d0 U285 ( .A(n221), .B(n232), .CI(n417), .CO(n418), .S(product[7]) );
  ad01d0 U286 ( .A(n233), .B(n246), .CI(n418), .CO(n419), .S(product[8]) );
  ad01d0 U287 ( .A(n247), .B(n262), .CI(n419), .CO(n420), .S(product[9]) );
  ad01d0 U288 ( .A(n263), .B(n280), .CI(n420), .CO(n421), .S(product[10]) );
  ad01d0 U289 ( .A(n281), .B(n300), .CI(n421), .CO(n422), .S(product[11]) );
  ad01d0 U290 ( .A(n301), .B(n320), .CI(n422), .CO(n423), .S(product[12]) );
  ad01d0 U291 ( .A(n321), .B(n338), .CI(n423), .CO(n424), .S(product[13]) );
  ad01d0 U292 ( .A(n339), .B(n354), .CI(n424), .CO(n425), .S(product[14]) );
  ad01d0 U293 ( .A(n355), .B(n368), .CI(n425), .CO(n426), .S(product[15]) );
  ad01d0 U296 ( .A(n398), .B(n391), .CI(n428), .CO(n429), .S(product[18]) );
  ad01d0 U297 ( .A(n404), .B(n399), .CI(n429), .CO(n430), .S(product[19]) );
  ad01d0 U298 ( .A(n408), .B(n405), .CI(n430), .CO(n431), .S(product[20]) );
  ad01d0 U299 ( .A(n410), .B(n409), .CI(n431), .CO(n432), .S(product[21]) );
  ad01d0 U300 ( .A(n191), .B(n411), .CI(n432), .CO(product[23]), .S(
        product[22]) );
  ad01d0 U304 ( .A(n369), .B(n380), .CI(n426), .CO(n427), .S(product[16]) );
  ad01d0 U305 ( .A(n390), .B(n381), .CI(n427), .CO(n428), .S(product[17]) );
  ah01d0 U306 ( .A(n50), .B(n61), .CO(n193), .S(n192) );
  ad01d0 U307 ( .A(n72), .B(n412), .CI(n192), .CO(n413), .S(product[2]) );
  inv0d1 U308 ( .I(a[0]), .ZN(n24) );
  inv0d1 U309 ( .I(a[5]), .ZN(n29) );
  inv0d1 U310 ( .I(a[4]), .ZN(n28) );
  inv0d1 U311 ( .I(a[2]), .ZN(n26) );
  inv0d1 U312 ( .I(a[3]), .ZN(n27) );
  inv0d1 U313 ( .I(a[1]), .ZN(n25) );
  inv0d1 U314 ( .I(b[0]), .ZN(n36) );
  inv0d1 U315 ( .I(b[1]), .ZN(n37) );
  inv0d1 U316 ( .I(b[3]), .ZN(n39) );
  inv0d1 U317 ( .I(b[4]), .ZN(n40) );
  inv0d1 U318 ( .I(b[2]), .ZN(n38) );
  inv0d1 U319 ( .I(a[6]), .ZN(n30) );
  inv0d1 U320 ( .I(a[7]), .ZN(n31) );
  inv0d1 U321 ( .I(a[8]), .ZN(n32) );
  inv0d1 U322 ( .I(a[9]), .ZN(n33) );
  inv0d1 U323 ( .I(a[10]), .ZN(n34) );
  inv0d1 U324 ( .I(b[8]), .ZN(n44) );
  inv0d1 U325 ( .I(b[10]), .ZN(n46) );
  inv0d1 U326 ( .I(b[9]), .ZN(n45) );
  inv0d1 U327 ( .I(b[11]), .ZN(n47) );
  inv0d1 U328 ( .I(b[5]), .ZN(n41) );
  inv0d1 U329 ( .I(b[6]), .ZN(n42) );
  inv0d1 U330 ( .I(b[7]), .ZN(n43) );
  inv0d1 U331 ( .I(a[11]), .ZN(n35) );
endmodule


module STACK_TOP ( reset_n, clk, PushEnbl, PopEnbl, PushDataIn, PopDataOut, 
        STACK_FULL, test_si, test_se, test_so );
  input [11:0] PushDataIn;
  output [11:0] PopDataOut;
  input reset_n, clk, PushEnbl, PopEnbl, test_si, test_se;
  output STACK_FULL, test_so;
  wire   n1, n2, n3, n4, n5, n6, n7, n10, n11, n12;
  wire   [0:2] TOS;

  STACK_FSM I_STACK_FSM ( .reset_n(reset_n), .clk(clk), .PushEnbl(n4), 
        .PopEnbl(PopEnbl), .TOS(TOS), .STACK_FULL(STACK_FULL), .test_se(
        test_se), .test_si(n10), .test_so(test_so) );
  STACK_MEM_0 I1_STACK_MEM ( .clk(clk), .PushEnbl(n5), .PopEnbl(PopEnbl), 
        .Stack_Full(STACK_FULL), .TOS({n3, n1, n2}), .PushDataIn(
        PushDataIn[3:0]), .PopDataOut(PopDataOut[3:0]), .test_se(test_se), 
        .test_si(test_si), .test_so(n12) );
  STACK_MEM_2 I2_STACK_MEM ( .clk(clk), .PushEnbl(n6), .PopEnbl(PopEnbl), 
        .Stack_Full(STACK_FULL), .TOS({n3, n1, n2}), .PushDataIn(
        PushDataIn[7:4]), .PopDataOut(PopDataOut[7:4]), .test_se(test_se), 
        .test_si(n12), .test_so(n11) );
  STACK_MEM_1 I3_STACK_MEM ( .clk(clk), .PushEnbl(n5), .PopEnbl(PopEnbl), 
        .Stack_Full(STACK_FULL), .TOS({n3, n1, n2}), .PushDataIn(
        PushDataIn[11:8]), .PopDataOut(PopDataOut[11:8]), .test_se(test_se), 
        .test_si(n11), .test_so(n10) );
  bufbd1 U1 ( .I(TOS[1]), .Z(n1) );
  bufbd1 U2 ( .I(TOS[2]), .Z(n2) );
  bufbd1 U3 ( .I(TOS[0]), .Z(n3) );
  inv0d1 U4 ( .I(n7), .ZN(n5) );
  inv0d1 U5 ( .I(n7), .ZN(n4) );
  inv0d1 U6 ( .I(n7), .ZN(n6) );
  inv0d1 U7 ( .I(PushEnbl), .ZN(n7) );
endmodule


module REG_FILE ( reset_n, clk, Addr_A, Addr_B, Addr_C, RegPort_C, Write_RegC, 
        RegPort_A, RegPort_B );
  input [6:0] Addr_A;
  input [6:0] Addr_B;
  input [6:0] Addr_C;
  input [15:0] RegPort_C;
  output [15:0] RegPort_A;
  output [15:0] RegPort_B;
  input reset_n, clk, Write_RegC;
  wire   we_n, SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192;

  ram16x128 REG_FILE_A_RAM ( .A1(Addr_C), .A2(Addr_A), .I1(RegPort_C), .O1({
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .O2({RegPort_A[15:8], SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120}), .CE1(clk), .CE2(clk), .OEB1(1'b1), .OEB2(
        1'b0), .CSB1(1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram16x128 REG_FILE_B_RAM ( .A1(Addr_C), .A2(Addr_B), .I1(RegPort_C), .O1({
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, 
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, 
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .O2({RegPort_B[15:8], SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144}), .CE1(clk), .CE2(clk), .OEB1(1'b1), .OEB2(
        1'b0), .CSB1(1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram16x128 REG_FILE_C_RAM ( .A1(Addr_C), .A2(Addr_A), .I1(RegPort_C), .O1({
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .O2({SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, RegPort_A[7:0]}), 
        .CE1(clk), .CE2(clk), .OEB1(1'b1), .OEB2(1'b0), .CSB1(1'b0), .CSB2(
        1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram16x128 REG_FILE_D_RAM ( .A1(Addr_C), .A2(Addr_B), .I1(RegPort_C), .O1({
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .O2({SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, RegPort_B[7:0]}), 
        .CE1(clk), .CE2(clk), .OEB1(1'b1), .OEB2(1'b0), .CSB1(1'b0), .CSB2(
        1'b0), .WEB1(we_n), .WEB2(1'b1) );
  inv0d1 U3 ( .I(Write_RegC), .ZN(we_n) );
endmodule


module PRGRM_CNT_TOP ( clk, reset_n, Crnt_Instrn, Zro_Flag, Carry_Flag, 
        Neg_Flag, Return_Addr, Current_State, PC, test_si, test_se );
  input [31:0] Crnt_Instrn;
  input [7:0] Return_Addr;
  output [2:0] Current_State;
  output [7:0] PC;
  input clk, reset_n, Zro_Flag, Carry_Flag, Neg_Flag, test_si, test_se;
  wire   Incrmnt_PC, Ld_Brnch_Addr, Ld_Rtn_Addr;

  PRGRM_FSM I_PRGRM_FSM ( .clk(clk), .reset_n(reset_n), .CurrentState(
        Current_State), .test_se(test_se), .test_si(PC[7]) );
  PRGRM_DECODE I_PRGRM_DECODE ( .Zro_Flag(Zro_Flag), .Carry_Flag(Carry_Flag), 
        .Neg_Flag(Neg_Flag), .CurrentState(Current_State), .Crnt_Instrn(
        Crnt_Instrn), .Incrmnt_PC(Incrmnt_PC), .Ld_Brnch_Addr(Ld_Brnch_Addr), 
        .Ld_Rtn_Addr(Ld_Rtn_Addr) );
  PRGRM_CNT I_PRGRM_CNT ( .reset_n(reset_n), .clk(clk), .Incrmnt_PC(Incrmnt_PC), .Ld_Brnch_Addr(Ld_Brnch_Addr), .Ld_Rtn_Addr(Ld_Rtn_Addr), .Imm_Addr(
        Crnt_Instrn[7:0]), .Return_Addr(Return_Addr), .PC(PC), .test_se(
        test_se), .test_si(test_si) );
endmodule


module INSTRN_LAT ( clk, Instrn, Latch_Instr, Crnt_Instrn_1, Crnt_Instrn_2, 
        test_se, test_si1, test_si2 );
  input [31:0] Instrn;
  output [31:0] Crnt_Instrn_1;
  output [31:0] Crnt_Instrn_2;
  input clk, Latch_Instr, test_se, test_si1, test_si2;
  wire   n64, n66, n67, n68, n69, n70, n71;

  senrq1 Crnt_Instrn_1_reg_10_ ( .D(Instrn[10]), .SD(Crnt_Instrn_1[9]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[10]) );
  senrq1 Crnt_Instrn_1_reg_14_ ( .D(Instrn[14]), .SD(Crnt_Instrn_1[13]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[14]) );
  senrq1 Crnt_Instrn_1_reg_13_ ( .D(Instrn[13]), .SD(Crnt_Instrn_1[12]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[13]) );
  senrq1 Crnt_Instrn_1_reg_12_ ( .D(Instrn[12]), .SD(Crnt_Instrn_1[11]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[12]) );
  senrq1 Crnt_Instrn_1_reg_11_ ( .D(Instrn[11]), .SD(Crnt_Instrn_1[10]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[11]) );
  senrq1 Crnt_Instrn_1_reg_8_ ( .D(Instrn[8]), .SD(Crnt_Instrn_1[7]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[8]) );
  senrq1 Crnt_Instrn_1_reg_7_ ( .D(Instrn[7]), .SD(Crnt_Instrn_1[6]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[7]) );
  senrq1 Crnt_Instrn_1_reg_15_ ( .D(Instrn[15]), .SD(Crnt_Instrn_1[14]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[15]) );
  senrq1 Crnt_Instrn_1_reg_9_ ( .D(Instrn[9]), .SD(Crnt_Instrn_1[8]), .ENN(n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[9]) );
  senrq1 Crnt_Instrn_2_reg_15_ ( .D(Instrn[15]), .SD(Crnt_Instrn_2[14]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[15]) );
  senrq1 Crnt_Instrn_2_reg_14_ ( .D(Instrn[14]), .SD(Crnt_Instrn_2[13]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[14]) );
  senrq1 Crnt_Instrn_2_reg_13_ ( .D(Instrn[13]), .SD(Crnt_Instrn_2[12]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[13]) );
  senrq1 Crnt_Instrn_2_reg_12_ ( .D(Instrn[12]), .SD(Crnt_Instrn_2[11]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[12]) );
  senrq1 Crnt_Instrn_2_reg_11_ ( .D(Instrn[11]), .SD(Crnt_Instrn_2[10]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[11]) );
  senrq1 Crnt_Instrn_2_reg_10_ ( .D(Instrn[10]), .SD(Crnt_Instrn_2[9]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[10]) );
  senrq1 Crnt_Instrn_2_reg_9_ ( .D(Instrn[9]), .SD(Crnt_Instrn_2[8]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[9]) );
  senrq1 Crnt_Instrn_2_reg_8_ ( .D(Instrn[8]), .SD(Crnt_Instrn_2[7]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[8]) );
  senrq1 Crnt_Instrn_1_reg_31_ ( .D(Instrn[31]), .SD(Crnt_Instrn_1[30]), .ENN(
        n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[31]) );
  senrq1 Crnt_Instrn_1_reg_30_ ( .D(Instrn[30]), .SD(Crnt_Instrn_1[29]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[30]) );
  senrq1 Crnt_Instrn_1_reg_23_ ( .D(Instrn[23]), .SD(Crnt_Instrn_1[22]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[23]) );
  senrq1 Crnt_Instrn_2_reg_7_ ( .D(Instrn[7]), .SD(Crnt_Instrn_2[6]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[7]) );
  senrq1 Crnt_Instrn_1_reg_29_ ( .D(Instrn[29]), .SD(Crnt_Instrn_1[28]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[29]) );
  senrq1 Crnt_Instrn_2_reg_6_ ( .D(Instrn[6]), .SD(Crnt_Instrn_2[5]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[6]) );
  senrq1 Crnt_Instrn_2_reg_5_ ( .D(Instrn[5]), .SD(Crnt_Instrn_2[4]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[5]) );
  senrq1 Crnt_Instrn_2_reg_4_ ( .D(Instrn[4]), .SD(Crnt_Instrn_2[3]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[4]) );
  senrq1 Crnt_Instrn_2_reg_3_ ( .D(Instrn[3]), .SD(Crnt_Instrn_2[2]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[3]) );
  senrq1 Crnt_Instrn_2_reg_2_ ( .D(Instrn[2]), .SD(Crnt_Instrn_2[1]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[2]) );
  senrq1 Crnt_Instrn_2_reg_1_ ( .D(Instrn[1]), .SD(Crnt_Instrn_2[0]), .ENN(n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[1]) );
  senrq1 Crnt_Instrn_2_reg_0_ ( .D(Instrn[0]), .SD(Crnt_Instrn_1[31]), .ENN(
        n68), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[0]) );
  senrq1 Crnt_Instrn_1_reg_6_ ( .D(Instrn[6]), .SD(Crnt_Instrn_1[5]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[6]) );
  senrq1 Crnt_Instrn_1_reg_5_ ( .D(Instrn[5]), .SD(Crnt_Instrn_1[4]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[5]) );
  senrq1 Crnt_Instrn_1_reg_4_ ( .D(Instrn[4]), .SD(Crnt_Instrn_1[3]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[4]) );
  senrq1 Crnt_Instrn_1_reg_3_ ( .D(Instrn[3]), .SD(test_si2), .ENN(n71), .SC(
        test_se), .CP(clk), .Q(Crnt_Instrn_1[3]) );
  senrq1 Crnt_Instrn_1_reg_2_ ( .D(Instrn[2]), .SD(Crnt_Instrn_1[1]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[2]) );
  senrq1 Crnt_Instrn_1_reg_22_ ( .D(Instrn[22]), .SD(Crnt_Instrn_1[21]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[22]) );
  senrq1 Crnt_Instrn_1_reg_21_ ( .D(Instrn[21]), .SD(Crnt_Instrn_1[20]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[21]) );
  senrq1 Crnt_Instrn_1_reg_20_ ( .D(Instrn[20]), .SD(Crnt_Instrn_1[19]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[20]) );
  senrq1 Crnt_Instrn_1_reg_19_ ( .D(Instrn[19]), .SD(Crnt_Instrn_1[18]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[19]) );
  senrq1 Crnt_Instrn_1_reg_18_ ( .D(Instrn[18]), .SD(Crnt_Instrn_1[17]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[18]) );
  senrq1 Crnt_Instrn_1_reg_17_ ( .D(Instrn[17]), .SD(Crnt_Instrn_1[16]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[17]) );
  senrq1 Crnt_Instrn_1_reg_16_ ( .D(Instrn[16]), .SD(Crnt_Instrn_1[15]), .ENN(
        n70), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[16]) );
  senrq1 Crnt_Instrn_1_reg_0_ ( .D(Instrn[0]), .SD(test_si1), .ENN(n71), .SC(
        test_se), .CP(clk), .Q(Crnt_Instrn_1[0]) );
  senrq1 Crnt_Instrn_1_reg_1_ ( .D(Instrn[1]), .SD(Crnt_Instrn_1[0]), .ENN(n71), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[1]) );
  senrq1 Crnt_Instrn_1_reg_25_ ( .D(Instrn[25]), .SD(Crnt_Instrn_1[24]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[25]) );
  senrq1 Crnt_Instrn_1_reg_24_ ( .D(Instrn[24]), .SD(Crnt_Instrn_1[23]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[24]) );
  senrq1 Crnt_Instrn_2_reg_26_ ( .D(Instrn[26]), .SD(Crnt_Instrn_2[25]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[26]) );
  senrq1 Crnt_Instrn_2_reg_29_ ( .D(Instrn[29]), .SD(Crnt_Instrn_2[28]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[29]) );
  senrq1 Crnt_Instrn_2_reg_27_ ( .D(Instrn[27]), .SD(Crnt_Instrn_2[26]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[27]) );
  senrq1 Crnt_Instrn_2_reg_24_ ( .D(Instrn[24]), .SD(Crnt_Instrn_2[23]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[24]) );
  senrq1 Crnt_Instrn_2_reg_21_ ( .D(Instrn[21]), .SD(Crnt_Instrn_2[20]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[21]) );
  senrq1 Crnt_Instrn_2_reg_19_ ( .D(Instrn[19]), .SD(Crnt_Instrn_2[18]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[19]) );
  senrq1 Crnt_Instrn_2_reg_18_ ( .D(Instrn[18]), .SD(Crnt_Instrn_2[17]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[18]) );
  senrq1 Crnt_Instrn_2_reg_20_ ( .D(Instrn[20]), .SD(Crnt_Instrn_2[19]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[20]) );
  senrq1 Crnt_Instrn_2_reg_23_ ( .D(Instrn[23]), .SD(Crnt_Instrn_2[22]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[23]) );
  senrq1 Crnt_Instrn_2_reg_22_ ( .D(Instrn[22]), .SD(Crnt_Instrn_2[21]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[22]) );
  senrq1 Crnt_Instrn_2_reg_16_ ( .D(Instrn[16]), .SD(Crnt_Instrn_2[15]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[16]) );
  senrq1 Crnt_Instrn_2_reg_17_ ( .D(Instrn[17]), .SD(Crnt_Instrn_2[16]), .ENN(
        n67), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[17]) );
  senrq1 Crnt_Instrn_1_reg_27_ ( .D(Instrn[27]), .SD(Crnt_Instrn_1[26]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[27]) );
  senrq1 Crnt_Instrn_2_reg_28_ ( .D(Instrn[28]), .SD(Crnt_Instrn_2[27]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[28]) );
  senrq1 Crnt_Instrn_1_reg_26_ ( .D(Instrn[26]), .SD(Crnt_Instrn_1[25]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[26]) );
  senrq1 Crnt_Instrn_1_reg_28_ ( .D(Instrn[28]), .SD(Crnt_Instrn_1[27]), .ENN(
        n69), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_1[28]) );
  senrq1 Crnt_Instrn_2_reg_25_ ( .D(Instrn[25]), .SD(Crnt_Instrn_2[24]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[25]) );
  senrq1 Crnt_Instrn_2_reg_31_ ( .D(Instrn[31]), .SD(Crnt_Instrn_2[30]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[31]) );
  senrq1 Crnt_Instrn_2_reg_30_ ( .D(Instrn[30]), .SD(Crnt_Instrn_2[29]), .ENN(
        n66), .SC(test_se), .CP(clk), .Q(Crnt_Instrn_2[30]) );
  bufbd1 U65 ( .I(n64), .Z(n70) );
  bufbd1 U67 ( .I(n64), .Z(n69) );
  bufbd1 U68 ( .I(n64), .Z(n68) );
  bufbd1 U69 ( .I(n64), .Z(n67) );
  bufbd1 U70 ( .I(n64), .Z(n66) );
  bufbd1 U71 ( .I(n64), .Z(n71) );
  inv0d1 U72 ( .I(Latch_Instr), .ZN(n64) );
endmodule


module DATA_PATH ( clk, reset_n, Reset_AluRegs, Rd_Oprnd_A, Rd_Oprnd_B, 
        UseData_Imm_Or_RegB, UseData_Imm_Or_ALU, Latch_Flags, ALU_Zro, ALU_Neg, 
        ALU_Carry, PSW_Zro, PSW_Neg, PSW_Carry, Crnt_Instrn, RegPort_A, 
        RegPort_B, Op_Result, Zro_Flag, Neg_Flag, Carry_Flag, Addr_A, Oprnd_A, 
        Oprnd_B, RegPort_C, test_se, test_si, test_so );
  input [31:0] Crnt_Instrn;
  input [15:0] RegPort_A;
  input [15:0] RegPort_B;
  input [15:0] Op_Result;
  output [6:0] Addr_A;
  output [15:0] Oprnd_A;
  output [15:0] Oprnd_B;
  output [15:0] RegPort_C;
  input clk, reset_n, Reset_AluRegs, Rd_Oprnd_A, Rd_Oprnd_B,
         UseData_Imm_Or_RegB, UseData_Imm_Or_ALU, Latch_Flags, ALU_Zro,
         ALU_Neg, ALU_Carry, PSW_Zro, PSW_Neg, PSW_Carry, test_se, test_si;
  output Zro_Flag, Neg_Flag, Carry_Flag, test_so;
  wire   N12, N14, N16, N18, N20, N22, N24, N26, N28, N30, N32, N34, N36, N38,
         N40, N41, N42, N94, N96, N98, N99, N100, N102, N104, N106, N108, N110,
         N112, N114, N116, N118, N120, N122, N124, PSWL_Neg, PSWL_Carry, n4,
         n21, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n1,
         n51;

  an02d1 U42 ( .A1(RegPort_A[15]), .A2(n45), .Z(N42) );
  an02d1 U43 ( .A1(RegPort_A[14]), .A2(n45), .Z(N40) );
  an02d1 U44 ( .A1(RegPort_A[13]), .A2(n45), .Z(N38) );
  an02d1 U45 ( .A1(RegPort_A[12]), .A2(n45), .Z(N36) );
  an02d1 U46 ( .A1(RegPort_A[11]), .A2(n45), .Z(N34) );
  an02d1 U47 ( .A1(RegPort_A[10]), .A2(n45), .Z(N32) );
  an02d1 U48 ( .A1(RegPort_A[9]), .A2(n45), .Z(N30) );
  an02d1 U49 ( .A1(RegPort_A[8]), .A2(n45), .Z(N28) );
  an02d1 U50 ( .A1(RegPort_A[7]), .A2(n45), .Z(N26) );
  an02d1 U51 ( .A1(RegPort_A[6]), .A2(n45), .Z(N24) );
  an02d1 U52 ( .A1(RegPort_A[5]), .A2(n45), .Z(N22) );
  an02d1 U53 ( .A1(RegPort_A[4]), .A2(n45), .Z(N20) );
  an02d1 U54 ( .A1(RegPort_A[3]), .A2(n45), .Z(N18) );
  an02d1 U55 ( .A1(RegPort_A[2]), .A2(n45), .Z(N16) );
  an02d1 U56 ( .A1(RegPort_A[1]), .A2(n45), .Z(N14) );
  an02d1 U57 ( .A1(RegPort_B[15]), .A2(n51), .Z(N124) );
  an02d1 U58 ( .A1(RegPort_B[14]), .A2(n51), .Z(N122) );
  an02d1 U59 ( .A1(RegPort_B[13]), .A2(n51), .Z(N120) );
  an02d1 U60 ( .A1(RegPort_A[0]), .A2(n45), .Z(N12) );
  an02d1 U61 ( .A1(RegPort_B[12]), .A2(n51), .Z(N118) );
  an02d1 U62 ( .A1(RegPort_B[11]), .A2(n51), .Z(N116) );
  an02d1 U63 ( .A1(RegPort_B[10]), .A2(n51), .Z(N114) );
  an02d1 U64 ( .A1(RegPort_B[9]), .A2(n51), .Z(N112) );
  an02d1 U65 ( .A1(RegPort_B[8]), .A2(n51), .Z(N110) );
  an02d1 U68 ( .A1(UseData_Imm_Or_RegB), .A2(n45), .Z(n44) );
  aor22d1 U73 ( .A1(test_so), .A2(n40), .B1(ALU_Zro), .B2(n41), .Z(Zro_Flag)
         );
  aor22d1 U74 ( .A1(Op_Result[9]), .A2(n42), .B1(n1), .B2(Crnt_Instrn[9]), .Z(
        RegPort_C[9]) );
  aor22d1 U75 ( .A1(Op_Result[8]), .A2(n42), .B1(Crnt_Instrn[8]), .B2(n1), .Z(
        RegPort_C[8]) );
  aor22d1 U76 ( .A1(Op_Result[7]), .A2(n42), .B1(Crnt_Instrn[7]), .B2(n1), .Z(
        RegPort_C[7]) );
  aor22d1 U77 ( .A1(Op_Result[6]), .A2(n42), .B1(Crnt_Instrn[6]), .B2(n1), .Z(
        RegPort_C[6]) );
  aor22d1 U78 ( .A1(Op_Result[5]), .A2(n42), .B1(Crnt_Instrn[5]), .B2(n1), .Z(
        RegPort_C[5]) );
  aor22d1 U79 ( .A1(Op_Result[4]), .A2(n42), .B1(Crnt_Instrn[4]), .B2(n1), .Z(
        RegPort_C[4]) );
  aor22d1 U80 ( .A1(Op_Result[3]), .A2(n42), .B1(Crnt_Instrn[3]), .B2(n1), .Z(
        RegPort_C[3]) );
  aor22d1 U81 ( .A1(Op_Result[2]), .A2(n42), .B1(Crnt_Instrn[2]), .B2(n1), .Z(
        RegPort_C[2]) );
  aor22d1 U82 ( .A1(Op_Result[1]), .A2(n42), .B1(Crnt_Instrn[1]), .B2(n1), .Z(
        RegPort_C[1]) );
  aor22d1 U83 ( .A1(Op_Result[15]), .A2(n42), .B1(Crnt_Instrn[15]), .B2(n1), 
        .Z(RegPort_C[15]) );
  aor22d1 U84 ( .A1(Op_Result[14]), .A2(n42), .B1(Crnt_Instrn[14]), .B2(n1), 
        .Z(RegPort_C[14]) );
  aor22d1 U85 ( .A1(Op_Result[13]), .A2(n42), .B1(Crnt_Instrn[13]), .B2(n1), 
        .Z(RegPort_C[13]) );
  aor22d1 U86 ( .A1(Op_Result[12]), .A2(n42), .B1(Crnt_Instrn[12]), .B2(n1), 
        .Z(RegPort_C[12]) );
  aor22d1 U87 ( .A1(Op_Result[11]), .A2(n42), .B1(Crnt_Instrn[11]), .B2(n1), 
        .Z(RegPort_C[11]) );
  aor22d1 U88 ( .A1(Op_Result[10]), .A2(n42), .B1(Crnt_Instrn[10]), .B2(n1), 
        .Z(RegPort_C[10]) );
  aor22d1 U89 ( .A1(Op_Result[0]), .A2(n42), .B1(Crnt_Instrn[0]), .B2(n1), .Z(
        RegPort_C[0]) );
  aor22d1 U91 ( .A1(RegPort_B[2]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[2]), 
        .Z(N98) );
  aor22d1 U92 ( .A1(RegPort_B[1]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[1]), 
        .Z(N96) );
  aor22d1 U93 ( .A1(RegPort_B[0]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[0]), 
        .Z(N94) );
  aor22d1 U94 ( .A1(RegPort_B[7]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[7]), 
        .Z(N108) );
  aor22d1 U95 ( .A1(RegPort_B[6]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[6]), 
        .Z(N106) );
  aor22d1 U96 ( .A1(RegPort_B[5]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[5]), 
        .Z(N104) );
  aor22d1 U97 ( .A1(RegPort_B[4]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[4]), 
        .Z(N102) );
  aor22d1 U98 ( .A1(RegPort_B[3]), .A2(n51), .B1(n44), .B2(Crnt_Instrn[3]), 
        .Z(N100) );
  nr02d0 U99 ( .A1(Reset_AluRegs), .A2(UseData_Imm_Or_RegB), .ZN(n43) );
  aor22d1 U100 ( .A1(PSWL_Carry), .A2(n40), .B1(ALU_Carry), .B2(n41), .Z(
        Carry_Flag) );
  nr04d0 U102 ( .A1(Crnt_Instrn[31]), .A2(Crnt_Instrn[30]), .A3(
        Crnt_Instrn[29]), .A4(Crnt_Instrn[28]), .ZN(n48) );
  nr02d0 U103 ( .A1(Crnt_Instrn[26]), .A2(Crnt_Instrn[25]), .ZN(n47) );
  aor22d1 U104 ( .A1(n49), .A2(Crnt_Instrn[6]), .B1(Crnt_Instrn[14]), .B2(n50), 
        .Z(Addr_A[6]) );
  aor22d1 U105 ( .A1(n49), .A2(Crnt_Instrn[5]), .B1(Crnt_Instrn[13]), .B2(n50), 
        .Z(Addr_A[5]) );
  aor22d1 U106 ( .A1(n49), .A2(Crnt_Instrn[4]), .B1(Crnt_Instrn[12]), .B2(n50), 
        .Z(Addr_A[4]) );
  aor22d1 U107 ( .A1(n49), .A2(Crnt_Instrn[3]), .B1(Crnt_Instrn[11]), .B2(n50), 
        .Z(Addr_A[3]) );
  aor22d1 U108 ( .A1(n49), .A2(Crnt_Instrn[2]), .B1(Crnt_Instrn[10]), .B2(n50), 
        .Z(Addr_A[2]) );
  aor22d1 U109 ( .A1(n49), .A2(Crnt_Instrn[1]), .B1(Crnt_Instrn[9]), .B2(n50), 
        .Z(Addr_A[1]) );
  aor22d1 U110 ( .A1(n49), .A2(Crnt_Instrn[0]), .B1(Crnt_Instrn[8]), .B2(n50), 
        .Z(Addr_A[0]) );
  nr03d0 U111 ( .A1(Crnt_Instrn[30]), .A2(Crnt_Instrn[31]), .A3(n46), .ZN(n49)
         );
  senrq1 Oprnd_B_reg_14_ ( .D(N122), .SD(Oprnd_B[13]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[14]) );
  senrq1 Oprnd_A_reg_15_ ( .D(N42), .SD(Oprnd_A[14]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[15]) );
  senrq1 Oprnd_B_reg_15_ ( .D(N124), .SD(Oprnd_B[14]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[15]) );
  senrq1 Oprnd_B_reg_13_ ( .D(N120), .SD(Oprnd_B[12]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[13]) );
  senrq1 Oprnd_B_reg_12_ ( .D(N118), .SD(Oprnd_B[11]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[12]) );
  senrq1 Oprnd_A_reg_13_ ( .D(N38), .SD(Oprnd_A[12]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[13]) );
  senrq1 Oprnd_A_reg_12_ ( .D(N36), .SD(Oprnd_A[11]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[12]) );
  secrq4 PSWL_Carry_reg ( .D(PSW_Carry), .SD(Oprnd_B[15]), .ENN(n4), .SC(
        test_se), .CP(clk), .CDN(reset_n), .Q(PSWL_Carry) );
  secrq4 PSWL_Zro_reg ( .D(PSW_Zro), .SD(PSWL_Neg), .ENN(n4), .SC(test_se), 
        .CP(clk), .CDN(reset_n), .Q(test_so) );
  secrq4 PSWL_Neg_reg ( .D(PSW_Neg), .SD(PSWL_Carry), .ENN(n4), .SC(test_se), 
        .CP(clk), .CDN(reset_n), .Q(PSWL_Neg) );
  senrq1 Oprnd_A_reg_10_ ( .D(N32), .SD(Oprnd_A[9]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[10]) );
  senrq1 Oprnd_A_reg_9_ ( .D(N30), .SD(Oprnd_A[8]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[9]) );
  senrq1 Oprnd_A_reg_8_ ( .D(N28), .SD(Oprnd_A[7]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[8]) );
  senrq1 Oprnd_B_reg_10_ ( .D(N114), .SD(Oprnd_B[9]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[10]) );
  senrq1 Oprnd_B_reg_9_ ( .D(N112), .SD(Oprnd_B[8]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[9]) );
  senrq1 Oprnd_B_reg_8_ ( .D(N110), .SD(Oprnd_B[7]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[8]) );
  senrq1 Oprnd_B_reg_11_ ( .D(N116), .SD(Oprnd_B[10]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[11]) );
  senrq1 Oprnd_A_reg_11_ ( .D(N34), .SD(Oprnd_A[10]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[11]) );
  senrq2 Oprnd_A_reg_0_ ( .D(N12), .SD(test_si), .ENN(n38), .SC(test_se), .CP(
        clk), .Q(Oprnd_A[0]) );
  senrq1 Oprnd_A_reg_5_ ( .D(N22), .SD(Oprnd_A[4]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[5]) );
  senrq1 Oprnd_A_reg_4_ ( .D(N20), .SD(Oprnd_A[3]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[4]) );
  senrq1 Oprnd_B_reg_7_ ( .D(N108), .SD(Oprnd_B[6]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[7]) );
  senrq1 Oprnd_B_reg_2_ ( .D(N98), .SD(Oprnd_B[1]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[2]) );
  senrq1 Oprnd_B_reg_6_ ( .D(N106), .SD(Oprnd_B[5]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[6]) );
  senrq1 Oprnd_A_reg_14_ ( .D(N40), .SD(Oprnd_A[13]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[14]) );
  senrq1 Oprnd_A_reg_7_ ( .D(N26), .SD(Oprnd_A[6]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[7]) );
  senrq1 Oprnd_A_reg_3_ ( .D(N18), .SD(Oprnd_A[2]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[3]) );
  senrq1 Oprnd_A_reg_1_ ( .D(N14), .SD(Oprnd_A[0]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[1]) );
  senrq1 Oprnd_A_reg_6_ ( .D(N24), .SD(Oprnd_A[5]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[6]) );
  senrq1 Oprnd_A_reg_2_ ( .D(N16), .SD(Oprnd_A[1]), .ENN(n38), .SC(test_se), 
        .CP(clk), .Q(Oprnd_A[2]) );
  senrq1 Oprnd_B_reg_5_ ( .D(N104), .SD(Oprnd_B[4]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[5]) );
  senrq1 Oprnd_B_reg_4_ ( .D(N102), .SD(Oprnd_B[3]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[4]) );
  senrq1 Oprnd_B_reg_3_ ( .D(N100), .SD(Oprnd_B[2]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[3]) );
  senrq1 Oprnd_B_reg_1_ ( .D(N96), .SD(Oprnd_B[0]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[1]) );
  senrq1 Oprnd_B_reg_0_ ( .D(N94), .SD(Oprnd_A[15]), .ENN(n21), .SC(test_se), 
        .CP(clk), .Q(Oprnd_B[0]) );
  inv0d1 U5 ( .I(Latch_Flags), .ZN(n4) );
  inv0d1 U22 ( .I(n41), .ZN(n40) );
  inv0d1 U39 ( .I(Reset_AluRegs), .ZN(n45) );
  inv0d1 U41 ( .I(n49), .ZN(n50) );
  inv0d1 U66 ( .I(N99), .ZN(n21) );
  nd12d0 U67 ( .A1(Rd_Oprnd_B), .A2(n45), .ZN(N99) );
  inv0d1 U69 ( .I(n1), .ZN(n42) );
  aor22d1 U70 ( .A1(PSWL_Neg), .A2(n40), .B1(ALU_Neg), .B2(n41), .Z(Neg_Flag)
         );
  nd04d0 U71 ( .A1(Crnt_Instrn[27]), .A2(n46), .A3(n47), .A4(n48), .ZN(n41) );
  inv0d1 U72 ( .I(Crnt_Instrn[24]), .ZN(n46) );
  inv0d1 U90 ( .I(N41), .ZN(n38) );
  nd12d0 U101 ( .A1(Rd_Oprnd_A), .A2(n45), .ZN(N41) );
  bufbd1 U112 ( .I(UseData_Imm_Or_ALU), .Z(n1) );
  bufbd1 U113 ( .I(n43), .Z(n51) );
endmodule


module CONTROL ( clk, reset_n, Crnt_Instrn, Current_State, Neg_Flag, 
        Carry_Flag, Zro_Flag, Latch_Instr, Rd_Oprnd_A, Rd_Oprnd_B, Latch_Flags, 
        Latch_Result, Write_RegC, UseData_Imm_Or_RegB, UseData_Imm_Or_ALU, 
        Reset_AluRegs, EndOfInstrn, PushEnbl, PopEnbl, OUT_VALID, test_se, 
        test_si );
  input [31:0] Crnt_Instrn;
  input [2:0] Current_State;
  input clk, reset_n, Neg_Flag, Carry_Flag, Zro_Flag, test_se, test_si;
  output Latch_Instr, Rd_Oprnd_A, Rd_Oprnd_B, Latch_Flags, Latch_Result,
         Write_RegC, UseData_Imm_Or_RegB, UseData_Imm_Or_ALU, Reset_AluRegs,
         EndOfInstrn, PushEnbl, PopEnbl, OUT_VALID;
  wire   Data_Imm_Or_RegB, Data_Imm_Or_ALU, N87, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31;

  an03d1 U6 ( .A1(n11), .A2(n12), .A3(Crnt_Instrn[28]), .Z(PushEnbl) );
  an02d1 U10 ( .A1(n22), .A2(n23), .Z(n16) );
  an04d1 U13 ( .A1(Crnt_Instrn[18]), .A2(Crnt_Instrn[19]), .A3(Crnt_Instrn[20]), .A4(Crnt_Instrn[21]), .Z(n20) );
  an02d1 U14 ( .A1(Crnt_Instrn[16]), .A2(n22), .Z(n18) );
  or04d1 U15 ( .A1(Crnt_Instrn[23]), .A2(Crnt_Instrn[22]), .A3(Crnt_Instrn[21]), .A4(Crnt_Instrn[20]), .Z(n25) );
  an02d1 U16 ( .A1(Crnt_Instrn[27]), .A2(n11), .Z(PopEnbl) );
  an03d1 U21 ( .A1(n8), .A2(n6), .A3(n27), .Z(n29) );
  nr02d0 U26 ( .A1(n5), .A2(n6), .ZN(Write_RegC) );
  nr03d0 U27 ( .A1(n7), .A2(Current_State[2]), .A3(Current_State[1]), .ZN(
        Reset_AluRegs) );
  nr02d0 U28 ( .A1(n5), .A2(n8), .ZN(Rd_Oprnd_B) );
  oan211d1 U29 ( .C1(Crnt_Instrn[30]), .C2(n9), .B(n10), .A(n8), .ZN(
        Rd_Oprnd_A) );
  aor22d1 U30 ( .A1(n13), .A2(n14), .B1(Crnt_Instrn[25]), .B2(n15), .Z(n12) );
  aor22d1 U31 ( .A1(n16), .A2(n17), .B1(n18), .B2(n19), .Z(n15) );
  aor222d1 U32 ( .A1(Zro_Flag), .A2(n18), .B1(n20), .B2(n21), .C1(Neg_Flag), 
        .C2(n16), .Z(n13) );
  nr04d0 U33 ( .A1(Crnt_Instrn[23]), .A2(Crnt_Instrn[22]), .A3(n23), .A4(n24), 
        .ZN(n21) );
  nr04d0 U34 ( .A1(Crnt_Instrn[18]), .A2(Crnt_Instrn[19]), .A3(Crnt_Instrn[17]), .A4(n25), .ZN(n22) );
  nr02d0 U35 ( .A1(n9), .A2(n26), .ZN(OUT_VALID) );
  nr02d0 U36 ( .A1(n5), .A2(n27), .ZN(Latch_Result) );
  nr02d0 U37 ( .A1(Crnt_Instrn[31]), .A2(Crnt_Instrn[30]), .ZN(n5) );
  nr02d0 U38 ( .A1(n10), .A2(n27), .ZN(Latch_Flags) );
  xn02d1 U39 ( .A1(Crnt_Instrn[30]), .A2(Crnt_Instrn[31]), .ZN(n10) );
  nr03d0 U40 ( .A1(n28), .A2(Crnt_Instrn[30]), .A3(n29), .ZN(Data_Imm_Or_RegB)
         );
  nr03d0 U41 ( .A1(n30), .A2(n29), .A3(n28), .ZN(Data_Imm_Or_ALU) );
  nd03d0 U42 ( .A1(Current_State[0]), .A2(n31), .A3(Current_State[1]), .ZN(n27) );
  nr03d0 U43 ( .A1(Current_State[0]), .A2(Current_State[1]), .A3(n31), .ZN(N87) );
  nd03d0 U44 ( .A1(n7), .A2(n31), .A3(Current_State[1]), .ZN(n8) );
  sdcrq1 UseData_Imm_Or_ALU_reg ( .D(Data_Imm_Or_ALU), .SD(EndOfInstrn), .SC(
        test_se), .CP(clk), .CDN(reset_n), .Q(UseData_Imm_Or_ALU) );
  sdcrq1 UseData_Imm_Or_RegB_reg ( .D(Data_Imm_Or_RegB), .SD(
        UseData_Imm_Or_ALU), .SC(test_se), .CP(clk), .CDN(reset_n), .Q(
        UseData_Imm_Or_RegB) );
  sdnrq1 EndOfInstrn_reg ( .D(N87), .SD(test_si), .SC(test_se), .CP(clk), .Q(
        EndOfInstrn) );
  inv0d0 U7 ( .I(Zro_Flag), .ZN(n19) );
  inv0d0 U8 ( .I(Neg_Flag), .ZN(n17) );
  inv0d0 U9 ( .I(Crnt_Instrn[24]), .ZN(n9) );
  inv0d0 U11 ( .I(Crnt_Instrn[25]), .ZN(n14) );
  inv0d0 U12 ( .I(Crnt_Instrn[30]), .ZN(n30) );
  inv0d0 U17 ( .I(Crnt_Instrn[31]), .ZN(n28) );
  inv0d1 U18 ( .I(n26), .ZN(n11) );
  nd12d0 U19 ( .A1(n27), .A2(n5), .ZN(n26) );
  inv0d1 U20 ( .I(N87), .ZN(n6) );
  inv0d1 U22 ( .I(Crnt_Instrn[17]), .ZN(n24) );
  inv0d1 U23 ( .I(Current_State[2]), .ZN(n31) );
  inv0d1 U24 ( .I(Current_State[0]), .ZN(n7) );
  inv0d1 U25 ( .I(Crnt_Instrn[16]), .ZN(n23) );
  bufbd1 U45 ( .I(Reset_AluRegs), .Z(Latch_Instr) );
endmodule


module ALU ( reset_n, clk, Oprnd_A, Oprnd_B, ALU_OP, Latch_Result, Latch_Flags, 
        Lachd_Result, Zro_Flag, Neg_Flag, Carry_Flag, test_se, test_si );
  input [15:0] Oprnd_A;
  input [15:0] Oprnd_B;
  input [5:0] ALU_OP;
  output [15:0] Lachd_Result;
  input reset_n, clk, Latch_Result, Latch_Flags, test_se, test_si;
  output Zro_Flag, Neg_Flag, Carry_Flag;
  wire   ALU_Zro, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, n17, n34, n69, n70, n74, n75, n83, n84, n99, n100, n105,
         n107, n108, n109, n113, n115, n116, n121, n123, n124, n125, n129,
         n131, n132, n133, n171, n172, n179, n180, n181, n187, n188, n189,
         n203, n204, n206, n208, n209, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n71, n72, n73, n76, n77,
         n78, n79, n80, n81, n82, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n101, n102, n103, n104, n106, n110, n111,
         n112, n114, n117, n118, n119, n120, n122, n126, n127, n128, n130,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n173, n174, n175, n176, n177, n178, n182,
         n183, n184, n185, n186, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n205, n207, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8;
  wire   [15:0] Result;

  nr02d0 U83 ( .A1(n57), .A2(n380), .ZN(Result[6]) );
  nr02d0 U84 ( .A1(n57), .A2(n379), .ZN(Result[5]) );
  nr02d0 U85 ( .A1(n57), .A2(n13), .ZN(Result[4]) );
  nr02d0 U86 ( .A1(n57), .A2(n14), .ZN(Result[3]) );
  nr02d0 U87 ( .A1(n57), .A2(n378), .ZN(Result[2]) );
  nr02d0 U88 ( .A1(n57), .A2(n377), .ZN(Result[1]) );
  nr02d0 U95 ( .A1(n57), .A2(n49), .ZN(Result[0]) );
  aor221d1 U102 ( .B1(n67), .B2(n383), .C1(n74), .C2(n385), .A(n75), .Z(n70)
         );
  aor22d1 U103 ( .A1(n67), .A2(n382), .B1(n54), .B2(n385), .Z(n69) );
  aor221d1 U109 ( .B1(n66), .B2(n383), .C1(n74), .C2(n386), .A(n75), .Z(n84)
         );
  aor22d1 U110 ( .A1(n66), .A2(n382), .B1(n54), .B2(n386), .Z(n83) );
  aor221d1 U123 ( .B1(n68), .B2(n383), .C1(n74), .C2(n384), .A(n75), .Z(n100)
         );
  aor22d1 U124 ( .A1(n68), .A2(n382), .B1(n54), .B2(n384), .Z(n99) );
  aor221d1 U130 ( .B1(n61), .B2(n383), .C1(n74), .C2(n105), .A(n75), .Z(n108)
         );
  aor22d1 U131 ( .A1(n61), .A2(n382), .B1(n54), .B2(n105), .Z(n107) );
  aor221d1 U137 ( .B1(n60), .B2(n383), .C1(n74), .C2(n113), .A(n75), .Z(n116)
         );
  aor22d1 U138 ( .A1(n8), .A2(n382), .B1(n54), .B2(n113), .Z(n115) );
  aor221d1 U144 ( .B1(n59), .B2(n383), .C1(n74), .C2(n121), .A(n75), .Z(n124)
         );
  aor22d1 U145 ( .A1(n59), .A2(n382), .B1(n54), .B2(n121), .Z(n123) );
  aor221d1 U151 ( .B1(n58), .B2(n383), .C1(n74), .C2(n129), .A(n75), .Z(n132)
         );
  aor22d1 U152 ( .A1(n58), .A2(n382), .B1(n54), .B2(n129), .Z(n131) );
  aor221d1 U186 ( .B1(n65), .B2(n383), .C1(n74), .C2(n387), .A(n75), .Z(n172)
         );
  aor22d1 U187 ( .A1(n65), .A2(n382), .B1(n54), .B2(n387), .Z(n171) );
  aor221d1 U193 ( .B1(n10), .B2(n383), .C1(n74), .C2(n388), .A(n75), .Z(n180)
         );
  aor22d1 U194 ( .A1(n10), .A2(n382), .B1(n54), .B2(n388), .Z(n179) );
  aor221d1 U200 ( .B1(n63), .B2(n383), .C1(n74), .C2(n389), .A(n75), .Z(n188)
         );
  aor22d1 U201 ( .A1(n63), .A2(n382), .B1(n54), .B2(n389), .Z(n187) );
  nr04d0 U209 ( .A1(ALU_OP[4]), .A2(ALU_OP[3]), .A3(n394), .A4(n208), .ZN(n206) );
  xn02d1 U210 ( .A1(n393), .A2(ALU_OP[0]), .ZN(n208) );
  aor221d1 U212 ( .B1(n62), .B2(n383), .C1(n74), .C2(n390), .A(n75), .Z(n204)
         );
  aor22d1 U214 ( .A1(n62), .A2(n382), .B1(n54), .B2(n390), .Z(n203) );
  nr03d0 U217 ( .A1(n391), .A2(ALU_OP[2]), .A3(n392), .ZN(n209) );
  ALU_DW01_sub_3 sub_89 ( .A({Oprnd_A[15:11], n68, n67, n66, n65, n10, n12, 
        n62, n61, n7, n59, n58}), .B(Oprnd_B), .CI(1'b0), .DIFF({N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113}), .CO(SYNOPSYS_UNCONNECTED_5) );
  ALU_DW01_sub_2 sub_1_root_sub_92 ( .A({Oprnd_A[15:11], n68, n67, n66, n65, 
        n64, n11, n62, n61, n7, n59, n58}), .B(Oprnd_B), .CI(1'b1), .DIFF({
        N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, 
        N148, N147, N146, N145}), .CO(SYNOPSYS_UNCONNECTED_6) );
  ALU_DW01_add_3 add_1_root_add_80_2 ( .A({Oprnd_A[15:11], n68, n67, n66, n65, 
        n9, n63, n62, n61, n60, n59, n58}), .B(Oprnd_B), .CI(1'b1), .SUM({N96, 
        N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, 
        N81}), .CO(SYNOPSYS_UNCONNECTED_7) );
  ALU_DW01_add_2 add_77 ( .A({Oprnd_A[15:11], n68, n67, n66, n65, n9, n11, n62, 
        n61, n8, n59, n58}), .B(Oprnd_B), .CI(1'b0), .SUM({N64, N63, N62, N61, 
        N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49}), .CO(
        SYNOPSYS_UNCONNECTED_8) );
  ALU_DW01_dec_1 sub_95 ( .A({Oprnd_A[15:11], n68, n67, n66, n65, n10, n63, 
        n62, n61, n60, n59, n58}), .SUM({N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161}) );
  ALU_DW01_inc_1 add_86 ( .A({Oprnd_A[15:11], n68, n67, n66, n65, n64, n12, 
        n62, n61, n8, n59, n58}), .SUM({N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97}) );
  secrq4 Zro_Flag_reg ( .D(ALU_Zro), .SD(Neg_Flag), .ENN(n17), .SC(test_se), 
        .CP(clk), .CDN(reset_n), .Q(Zro_Flag) );
  senrq1 Lachd_Result_reg_15_ ( .D(n381), .SD(Lachd_Result[14]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[15]) );
  senrq1 Lachd_Result_reg_14_ ( .D(Result[14]), .SD(Lachd_Result[13]), .ENN(
        n34), .SC(test_se), .CP(clk), .Q(Lachd_Result[14]) );
  senrq1 Lachd_Result_reg_13_ ( .D(Result[13]), .SD(Lachd_Result[12]), .ENN(
        n34), .SC(test_se), .CP(clk), .Q(Lachd_Result[13]) );
  senrq1 Lachd_Result_reg_12_ ( .D(Result[12]), .SD(Lachd_Result[11]), .ENN(
        n34), .SC(test_se), .CP(clk), .Q(Lachd_Result[12]) );
  senrq1 Lachd_Result_reg_11_ ( .D(Result[11]), .SD(Lachd_Result[10]), .ENN(
        n34), .SC(test_se), .CP(clk), .Q(Lachd_Result[11]) );
  senrq1 Lachd_Result_reg_10_ ( .D(Result[10]), .SD(Lachd_Result[9]), .ENN(n34), .SC(test_se), .CP(clk), .Q(Lachd_Result[10]) );
  senrq1 Lachd_Result_reg_9_ ( .D(Result[9]), .SD(Lachd_Result[8]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[9]) );
  senrq1 Lachd_Result_reg_8_ ( .D(Result[8]), .SD(Lachd_Result[7]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[8]) );
  senrq1 Lachd_Result_reg_7_ ( .D(Result[7]), .SD(Lachd_Result[6]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[7]) );
  senrq1 Lachd_Result_reg_6_ ( .D(Result[6]), .SD(Lachd_Result[5]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[6]) );
  senrq1 Lachd_Result_reg_5_ ( .D(Result[5]), .SD(Lachd_Result[4]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[5]) );
  senrq1 Lachd_Result_reg_4_ ( .D(Result[4]), .SD(Lachd_Result[3]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[4]) );
  senrq1 Lachd_Result_reg_3_ ( .D(Result[3]), .SD(Lachd_Result[2]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[3]) );
  senrq1 Lachd_Result_reg_2_ ( .D(Result[2]), .SD(Lachd_Result[1]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[2]) );
  senrq1 Lachd_Result_reg_1_ ( .D(Result[1]), .SD(Lachd_Result[0]), .ENN(n34), 
        .SC(test_se), .CP(clk), .Q(Lachd_Result[1]) );
  senrq1 Lachd_Result_reg_0_ ( .D(Result[0]), .SD(test_si), .ENN(n34), .SC(
        test_se), .CP(clk), .Q(Lachd_Result[0]) );
  secrq4 Neg_Flag_reg ( .D(n381), .SD(Lachd_Result[15]), .ENN(n17), .SC(
        test_se), .CP(clk), .CDN(reset_n), .Q(Neg_Flag) );
  inv0d1 U4 ( .I(1'b1), .ZN(Carry_Flag) );
  bufbd4 U6 ( .I(Oprnd_A[0]), .Z(n58) );
  bufbd1 U7 ( .I(Oprnd_A[2]), .Z(n7) );
  bufbd2 U8 ( .I(Oprnd_A[4]), .Z(n62) );
  bufbd1 U26 ( .I(Oprnd_A[2]), .Z(n60) );
  nd12d0 U28 ( .A1(n342), .A2(N146), .ZN(n110) );
  nd12d0 U29 ( .A1(n342), .A2(N147), .ZN(n138) );
  nd12d0 U30 ( .A1(n342), .A2(N148), .ZN(n192) );
  nd12d0 U31 ( .A1(n342), .A2(N149), .ZN(n173) );
  nd12d0 U32 ( .A1(n342), .A2(N150), .ZN(n212) );
  nd12d0 U33 ( .A1(n342), .A2(N151), .ZN(n225) );
  nd12d0 U34 ( .A1(n342), .A2(N152), .ZN(n315) );
  nd12d0 U35 ( .A1(n342), .A2(N153), .ZN(n303) );
  nd12d0 U36 ( .A1(n342), .A2(N154), .ZN(n327) );
  nd12d0 U37 ( .A1(n342), .A2(N155), .ZN(n343) );
  an02d1 U38 ( .A1(n360), .A2(n362), .Z(n3) );
  or02d1 U39 ( .A1(n245), .A2(n244), .Z(n4) );
  an02d1 U40 ( .A1(n359), .A2(n3), .Z(n5) );
  an02d1 U41 ( .A1(n203), .A2(Oprnd_B[4]), .Z(n6) );
  bufbd1 U42 ( .I(Oprnd_A[2]), .Z(n8) );
  an03d1 U43 ( .A1(n249), .A2(n248), .A3(n56), .Z(n372) );
  bufbd1 U44 ( .I(Oprnd_A[6]), .Z(n10) );
  bufbd1 U45 ( .I(Oprnd_A[6]), .Z(n64) );
  bufbd1 U46 ( .I(Oprnd_A[6]), .Z(n9) );
  nr03d0 U47 ( .A1(n247), .A2(n246), .A3(n4), .ZN(n248) );
  nd02d1 U48 ( .A1(n361), .A2(n5), .ZN(n363) );
  bufbd2 U49 ( .I(Oprnd_A[1]), .Z(n59) );
  bufbd2 U50 ( .I(Oprnd_A[7]), .Z(n65) );
  bufbd2 U51 ( .I(Oprnd_A[3]), .Z(n61) );
  bufbd1 U52 ( .I(Oprnd_A[5]), .Z(n12) );
  bufbd1 U53 ( .I(Oprnd_A[5]), .Z(n11) );
  bufbd1 U54 ( .I(Oprnd_A[5]), .Z(n63) );
  an02d1 U55 ( .A1(n170), .A2(n49), .Z(n361) );
  an04d1 U56 ( .A1(n372), .A2(n371), .A3(n358), .A4(n357), .Z(n359) );
  bufbd2 U57 ( .I(Oprnd_A[8]), .Z(n66) );
  bufbd1 U58 ( .I(Oprnd_A[9]), .Z(n67) );
  nd12d1 U59 ( .A1(n57), .A2(n363), .ZN(ALU_Zro) );
  nd12d1 U60 ( .A1(n104), .A2(n103), .ZN(n151) );
  nd12d0 U61 ( .A1(n98), .A2(n97), .ZN(n101) );
  nd12d0 U62 ( .A1(n342), .A2(N160), .ZN(n81) );
  nd12d0 U63 ( .A1(n337), .A2(N128), .ZN(n80) );
  nd12d0 U64 ( .A1(n346), .A2(N96), .ZN(n76) );
  nd12d0 U65 ( .A1(n338), .A2(N64), .ZN(n77) );
  an03d1 U66 ( .A1(n191), .A2(n190), .A3(n186), .Z(n13) );
  inv0d0 U67 ( .I(n348), .ZN(n93) );
  inv0d0 U68 ( .I(n364), .ZN(n365) );
  inv0d0 U69 ( .I(n366), .ZN(n367) );
  inv0d0 U70 ( .I(n368), .ZN(n369) );
  inv0d0 U71 ( .I(n375), .ZN(n379) );
  inv0d0 U72 ( .I(n376), .ZN(n380) );
  an03d1 U73 ( .A1(n211), .A2(n210), .A3(n207), .Z(n14) );
  an04d1 U74 ( .A1(n300), .A2(n299), .A3(n298), .A4(n297), .Z(n15) );
  an02d1 U75 ( .A1(n324), .A2(n323), .Z(n36) );
  inv0d0 U76 ( .I(n66), .ZN(n386) );
  inv0d0 U77 ( .I(n67), .ZN(n385) );
  inv0d0 U78 ( .I(n58), .ZN(n129) );
  inv0d0 U79 ( .I(n60), .ZN(n113) );
  inv0d0 U80 ( .I(n59), .ZN(n121) );
  inv0d0 U81 ( .I(n61), .ZN(n105) );
  inv0d0 U82 ( .I(n64), .ZN(n388) );
  inv0d0 U89 ( .I(n62), .ZN(n390) );
  inv0d0 U90 ( .I(n65), .ZN(n387) );
  inv0d0 U91 ( .I(n12), .ZN(n389) );
  inv0d1 U92 ( .I(n38), .ZN(n75) );
  nd02d0 U93 ( .A1(n91), .A2(ALU_OP[2]), .ZN(n85) );
  nd12d0 U94 ( .A1(Oprnd_B[2]), .A2(n116), .ZN(n142) );
  nd02d0 U96 ( .A1(n115), .A2(Oprnd_B[2]), .ZN(n143) );
  nd02d0 U97 ( .A1(ALU_OP[2]), .A2(ALU_OP[4]), .ZN(n88) );
  nd12d0 U98 ( .A1(Oprnd_B[4]), .A2(n204), .ZN(n178) );
  nd02d0 U99 ( .A1(n179), .A2(Oprnd_B[6]), .ZN(n230) );
  nd02d0 U100 ( .A1(n131), .A2(Oprnd_B[0]), .ZN(n162) );
  nd02d1 U101 ( .A1(n107), .A2(Oprnd_B[3]), .ZN(n198) );
  nd02d1 U104 ( .A1(n123), .A2(Oprnd_B[1]), .ZN(n120) );
  an03d1 U105 ( .A1(ALU_OP[1]), .A2(n392), .A3(n391), .Z(n37) );
  inv0d0 U106 ( .I(Oprnd_B[6]), .ZN(n181) );
  inv0d0 U107 ( .I(Oprnd_B[0]), .ZN(n133) );
  or03d1 U108 ( .A1(n393), .A2(n391), .A3(n392), .Z(n38) );
  nd02d1 U111 ( .A1(n39), .A2(n315), .ZN(n316) );
  nd02d1 U112 ( .A1(N104), .A2(n341), .ZN(n39) );
  nd02d1 U113 ( .A1(n40), .A2(n303), .ZN(n304) );
  nd02d1 U114 ( .A1(N105), .A2(n341), .ZN(n40) );
  nd02d1 U115 ( .A1(n41), .A2(n343), .ZN(n344) );
  nd02d1 U116 ( .A1(N107), .A2(n341), .ZN(n41) );
  nd02d1 U117 ( .A1(n42), .A2(n327), .ZN(n328) );
  nd02d1 U118 ( .A1(N106), .A2(n341), .ZN(n42) );
  inv0d1 U119 ( .I(n292), .ZN(n341) );
  nd12d0 U120 ( .A1(n338), .A2(N51), .ZN(n137) );
  nd12d0 U121 ( .A1(n346), .A2(N83), .ZN(n136) );
  nd02d1 U122 ( .A1(n43), .A2(n192), .ZN(n193) );
  nd02d1 U125 ( .A1(N100), .A2(n341), .ZN(n43) );
  nd02d1 U126 ( .A1(n44), .A2(n173), .ZN(n174) );
  nd02d1 U127 ( .A1(N101), .A2(n341), .ZN(n44) );
  nd02d1 U128 ( .A1(n45), .A2(n225), .ZN(n226) );
  nd02d1 U129 ( .A1(N103), .A2(n341), .ZN(n45) );
  nd02d1 U132 ( .A1(n46), .A2(n212), .ZN(n213) );
  nd02d1 U133 ( .A1(N102), .A2(n341), .ZN(n46) );
  nd02d1 U134 ( .A1(n47), .A2(n138), .ZN(n139) );
  nd02d1 U135 ( .A1(N99), .A2(n341), .ZN(n47) );
  nd12d0 U136 ( .A1(n338), .A2(N52), .ZN(n196) );
  nd12d0 U139 ( .A1(n346), .A2(N84), .ZN(n195) );
  an02d1 U140 ( .A1(n110), .A2(n48), .Z(n118) );
  nd02d1 U141 ( .A1(N98), .A2(n341), .ZN(n48) );
  nd12d0 U142 ( .A1(n342), .A2(N145), .ZN(n154) );
  inv0d1 U143 ( .I(Latch_Flags), .ZN(n17) );
  an12d1 U146 ( .A2(N159), .A1(n342), .Z(n242) );
  an12d1 U147 ( .A2(N157), .A1(n342), .Z(n272) );
  an12d1 U148 ( .A2(N158), .A1(n342), .Z(n256) );
  an12d1 U149 ( .A2(N93), .A1(n346), .Z(n278) );
  an12d1 U150 ( .A2(N94), .A1(n346), .Z(n262) );
  an12d1 U153 ( .A2(N63), .A1(n338), .Z(n247) );
  an12d1 U154 ( .A2(N127), .A1(n337), .Z(n243) );
  an12d1 U155 ( .A2(N125), .A1(n337), .Z(n273) );
  an12d1 U156 ( .A2(N126), .A1(n337), .Z(n257) );
  nd12d0 U157 ( .A1(n347), .A2(N171), .ZN(n352) );
  nd12d0 U158 ( .A1(n347), .A2(N170), .ZN(n333) );
  nd12d0 U159 ( .A1(n347), .A2(N169), .ZN(n309) );
  nd12d0 U160 ( .A1(n57), .A2(n151), .ZN(n106) );
  nd12d0 U161 ( .A1(n346), .A2(N89), .ZN(n310) );
  nd12d0 U162 ( .A1(n346), .A2(N92), .ZN(n299) );
  nd12d0 U163 ( .A1(n338), .A2(N60), .ZN(n300) );
  nd12d0 U164 ( .A1(n292), .A2(N111), .ZN(n250) );
  nd12d0 U165 ( .A1(n346), .A2(N91), .ZN(n353) );
  nd12d0 U166 ( .A1(n346), .A2(N90), .ZN(n334) );
  nd12d0 U167 ( .A1(n346), .A2(N88), .ZN(n322) );
  nd12d0 U168 ( .A1(n364), .A2(n36), .ZN(n356) );
  nd12d0 U169 ( .A1(n342), .A2(N156), .ZN(n287) );
  nd12d0 U170 ( .A1(n337), .A2(N124), .ZN(n286) );
  nd12d0 U171 ( .A1(n338), .A2(N56), .ZN(n313) );
  nd12d0 U172 ( .A1(n337), .A2(N120), .ZN(n314) );
  nd12d0 U173 ( .A1(n337), .A2(N121), .ZN(n302) );
  nd12d0 U174 ( .A1(n338), .A2(N57), .ZN(n301) );
  nd12d0 U175 ( .A1(n337), .A2(N123), .ZN(n340) );
  nd12d0 U176 ( .A1(n338), .A2(N59), .ZN(n339) );
  nd12d0 U177 ( .A1(n337), .A2(N122), .ZN(n326) );
  nd12d0 U178 ( .A1(n338), .A2(N58), .ZN(n325) );
  inv0d1 U179 ( .I(N62), .ZN(n258) );
  inv0d1 U180 ( .I(N61), .ZN(n274) );
  nd02d1 U181 ( .A1(n78), .A2(n37), .ZN(n347) );
  nd02d1 U182 ( .A1(n55), .A2(n37), .ZN(n292) );
  an02d1 U183 ( .A1(n209), .A2(n394), .Z(n74) );
  nd03d0 U184 ( .A1(n393), .A2(n79), .A3(n91), .ZN(n338) );
  nd02d1 U185 ( .A1(n78), .A2(n79), .ZN(n342) );
  nd02d1 U188 ( .A1(n55), .A2(n79), .ZN(n346) );
  nd12d0 U189 ( .A1(n347), .A2(N164), .ZN(n200) );
  nd12d0 U190 ( .A1(n105), .A2(n348), .ZN(n201) );
  nd12d0 U191 ( .A1(n163), .A2(n182), .ZN(n165) );
  nd12d0 U192 ( .A1(n129), .A2(n348), .ZN(n166) );
  nd12d0 U195 ( .A1(n347), .A2(N163), .ZN(n145) );
  nd12d0 U196 ( .A1(n113), .A2(n348), .ZN(n146) );
  nd12d0 U197 ( .A1(n347), .A2(N162), .ZN(n126) );
  nd12d0 U198 ( .A1(n121), .A2(n348), .ZN(n127) );
  nd12d0 U199 ( .A1(n135), .A2(n134), .ZN(n373) );
  nd12d0 U202 ( .A1(n337), .A2(N114), .ZN(n117) );
  nr02d0 U203 ( .A1(n169), .A2(n50), .ZN(n49) );
  or02d1 U204 ( .A1(n168), .A2(n167), .Z(n50) );
  nd12d0 U205 ( .A1(n346), .A2(N87), .ZN(n228) );
  nd12d0 U206 ( .A1(n346), .A2(N86), .ZN(n215) );
  nd12d0 U207 ( .A1(n346), .A2(N85), .ZN(n176) );
  nd12d0 U208 ( .A1(n338), .A2(N55), .ZN(n229) );
  nd12d0 U211 ( .A1(n338), .A2(N54), .ZN(n216) );
  nd12d0 U213 ( .A1(n338), .A2(N53), .ZN(n177) );
  mx02d0 U215 ( .I0(n53), .I1(n348), .S(n64), .Z(n232) );
  nd12d0 U216 ( .A1(n347), .A2(N168), .ZN(n321) );
  mx02d0 U218 ( .I0(n53), .I1(n348), .S(n62), .Z(n185) );
  nd12d0 U219 ( .A1(n337), .A2(N113), .ZN(n159) );
  an02d1 U220 ( .A1(n181), .A2(n180), .Z(n51) );
  an02d1 U221 ( .A1(n189), .A2(n188), .Z(n52) );
  inv0d1 U222 ( .I(n68), .ZN(n384) );
  nd12d0 U223 ( .A1(n346), .A2(N82), .ZN(n111) );
  nd12d0 U224 ( .A1(n338), .A2(N50), .ZN(n112) );
  inv0d1 U225 ( .I(Latch_Result), .ZN(n34) );
  nd12d0 U226 ( .A1(n206), .A2(n92), .ZN(n348) );
  nd12d0 U227 ( .A1(n91), .A2(n90), .ZN(n92) );
  mx02d0 U228 ( .I0(n383), .I1(n382), .S(Oprnd_B[11]), .Z(n289) );
  inv0d1 U229 ( .I(ALU_OP[2]), .ZN(n393) );
  mx02d0 U230 ( .I0(n172), .I1(n171), .S(Oprnd_B[7]), .Z(n319) );
  mx02d0 U231 ( .I0(n53), .I1(n348), .S(n65), .Z(n318) );
  mx02d0 U232 ( .I0(n84), .I1(n83), .S(Oprnd_B[8]), .Z(n307) );
  mx02d0 U233 ( .I0(n53), .I1(n348), .S(n66), .Z(n306) );
  mx02d0 U234 ( .I0(n100), .I1(n99), .S(Oprnd_B[10]), .Z(n350) );
  mx02d0 U235 ( .I0(n53), .I1(n348), .S(n68), .Z(n349) );
  mx02d0 U236 ( .I0(n70), .I1(n69), .S(Oprnd_B[9]), .Z(n331) );
  mx02d0 U237 ( .I0(n53), .I1(n348), .S(n67), .Z(n330) );
  inv0d1 U238 ( .I(ALU_OP[4]), .ZN(n391) );
  mx02d0 U239 ( .I0(n271), .I1(n270), .S(Oprnd_A[12]), .Z(n283) );
  nd02d1 U240 ( .A1(n341), .A2(N109), .ZN(n282) );
  mx02d0 U241 ( .I0(n255), .I1(n254), .S(Oprnd_A[13]), .Z(n267) );
  nd02d1 U242 ( .A1(n341), .A2(N110), .ZN(n266) );
  inv0d1 U243 ( .I(ALU_OP[3]), .ZN(n392) );
  bufbd1 U244 ( .I(Oprnd_A[10]), .Z(n68) );
  nd12d0 U245 ( .A1(n292), .A2(N112), .ZN(n97) );
  nd12d0 U246 ( .A1(n292), .A2(N108), .ZN(n293) );
  mx02d0 U247 ( .I0(n291), .I1(n290), .S(Oprnd_A[11]), .Z(n294) );
  nd12d0 U248 ( .A1(n89), .A2(n38), .ZN(n90) );
  nd12d0 U249 ( .A1(Oprnd_B[15]), .A2(n75), .ZN(n71) );
  nd12d0 U250 ( .A1(n347), .A2(N176), .ZN(n72) );
  an12d1 U251 ( .A2(N95), .A1(n346), .Z(n246) );
  inv0d1 U252 ( .I(N173), .ZN(n275) );
  inv0d1 U253 ( .I(N174), .ZN(n259) );
  an12d1 U254 ( .A2(N175), .A1(n347), .Z(n245) );
  an03d1 U255 ( .A1(ALU_OP[4]), .A2(ALU_OP[3]), .A3(ALU_OP[1]), .Z(n53) );
  an03d1 U256 ( .A1(ALU_OP[1]), .A2(ALU_OP[4]), .A3(n392), .Z(n54) );
  nr03d0 U257 ( .A1(n85), .A2(ALU_OP[3]), .A3(n391), .ZN(n383) );
  nr02d0 U258 ( .A1(n87), .A2(n91), .ZN(n382) );
  mx02d0 U259 ( .I0(n74), .I1(n54), .S(Oprnd_B[12]), .Z(n268) );
  mx02d0 U260 ( .I0(n74), .I1(n54), .S(Oprnd_B[13]), .Z(n252) );
  nd03d0 U261 ( .A1(ALU_OP[0]), .A2(ALU_OP[2]), .A3(n79), .ZN(n337) );
  an12d1 U262 ( .A2(n75), .A1(Oprnd_B[14]), .Z(n244) );
  mx02d0 U263 ( .I0(n383), .I1(n382), .S(Oprnd_B[12]), .Z(n269) );
  mx02d0 U264 ( .I0(n383), .I1(n382), .S(Oprnd_B[13]), .Z(n253) );
  an02d1 U265 ( .A1(ALU_OP[0]), .A2(n393), .Z(n55) );
  mx02d0 U266 ( .I0(n74), .I1(n54), .S(Oprnd_B[14]), .Z(n238) );
  nd12d0 U267 ( .A1(Oprnd_B[11]), .A2(n75), .ZN(n284) );
  nd02d1 U268 ( .A1(n133), .A2(n132), .ZN(n161) );
  nd12d0 U269 ( .A1(n347), .A2(N172), .ZN(n285) );
  mx02d0 U270 ( .I0(n383), .I1(n382), .S(Oprnd_B[14]), .Z(n239) );
  mx02d0 U271 ( .I0(n383), .I1(n382), .S(Oprnd_B[15]), .Z(n94) );
  mx02d0 U272 ( .I0(n96), .I1(n95), .S(Oprnd_A[15]), .Z(n98) );
  nd12d0 U273 ( .A1(n53), .A2(n82), .ZN(n96) );
  nd12d0 U274 ( .A1(n94), .A2(n93), .ZN(n95) );
  nd12d0 U275 ( .A1(n347), .A2(N167), .ZN(n231) );
  nd12d0 U276 ( .A1(n347), .A2(N166), .ZN(n218) );
  nd02d1 U277 ( .A1(n187), .A2(Oprnd_B[5]), .ZN(n217) );
  nd02d1 U278 ( .A1(n109), .A2(n108), .ZN(n197) );
  nd02d1 U279 ( .A1(n125), .A2(n124), .ZN(n119) );
  nd12d0 U280 ( .A1(n346), .A2(N81), .ZN(n156) );
  bufbd1 U281 ( .I(ALU_OP[5]), .Z(n57) );
  inv0d1 U282 ( .I(Oprnd_B[3]), .ZN(n109) );
  inv0d1 U283 ( .I(Oprnd_B[1]), .ZN(n125) );
  inv0d1 U284 ( .I(Oprnd_B[5]), .ZN(n189) );
  an02d1 U285 ( .A1(n250), .A2(n251), .Z(n56) );
  mx02d0 U286 ( .I0(n241), .I1(n240), .S(Oprnd_A[14]), .Z(n251) );
  mx02d0 U287 ( .I0(n53), .I1(n348), .S(n12), .Z(n219) );
  nr03d0 U288 ( .A1(ALU_OP[4]), .A2(ALU_OP[3]), .A3(ALU_OP[1]), .ZN(n79) );
  inv0d1 U289 ( .I(ALU_OP[0]), .ZN(n91) );
  inv0d1 U290 ( .I(n85), .ZN(n78) );
  an02d1 U291 ( .A1(n72), .A2(n71), .Z(n73) );
  nd03d0 U292 ( .A1(n77), .A2(n76), .A3(n73), .ZN(n104) );
  nd02d1 U293 ( .A1(n81), .A2(n80), .ZN(n102) );
  mi02d0 U294 ( .I0(n74), .I1(n54), .S(Oprnd_B[15]), .ZN(n82) );
  nr03d0 U295 ( .A1(ALU_OP[2]), .A2(ALU_OP[3]), .A3(n391), .ZN(n86) );
  nr02d0 U296 ( .A1(n209), .A2(n86), .ZN(n87) );
  nr02d0 U297 ( .A1(n88), .A2(ALU_OP[3]), .ZN(n89) );
  nr02d0 U298 ( .A1(n102), .A2(n101), .ZN(n103) );
  inv0d1 U299 ( .I(n106), .ZN(n381) );
  an02d1 U300 ( .A1(n112), .A2(n111), .Z(n114) );
  nd03d0 U301 ( .A1(n118), .A2(n117), .A3(n114), .ZN(n135) );
  nd02d1 U302 ( .A1(n120), .A2(n119), .ZN(n130) );
  nd02d1 U303 ( .A1(n121), .A2(n53), .ZN(n122) );
  nd03d0 U304 ( .A1(n127), .A2(n126), .A3(n122), .ZN(n128) );
  nr02d0 U305 ( .A1(n130), .A2(n128), .ZN(n134) );
  nd02d1 U306 ( .A1(n137), .A2(n136), .ZN(n141) );
  inv0d1 U307 ( .I(n337), .ZN(n224) );
  an02d1 U308 ( .A1(N115), .A2(n224), .Z(n140) );
  nr03d0 U309 ( .A1(n141), .A2(n140), .A3(n139), .ZN(n150) );
  nd02d1 U310 ( .A1(n143), .A2(n142), .ZN(n148) );
  nd02d1 U311 ( .A1(n113), .A2(n53), .ZN(n144) );
  nd03d0 U312 ( .A1(n146), .A2(n145), .A3(n144), .ZN(n147) );
  nr02d0 U313 ( .A1(n148), .A2(n147), .ZN(n149) );
  nd02d1 U314 ( .A1(n150), .A2(n149), .ZN(n374) );
  nr02d0 U315 ( .A1(n373), .A2(n374), .ZN(n362) );
  inv0d1 U316 ( .I(n151), .ZN(n170) );
  inv0d1 U317 ( .I(N97), .ZN(n152) );
  nr02d0 U318 ( .A1(n292), .A2(n152), .ZN(n153) );
  an12d1 U319 ( .A2(n154), .A1(n153), .Z(n160) );
  inv0d1 U320 ( .I(n338), .ZN(n155) );
  nd02d1 U321 ( .A1(N49), .A2(n155), .ZN(n157) );
  an02d1 U322 ( .A1(n157), .A2(n156), .Z(n158) );
  nd03d0 U323 ( .A1(n160), .A2(n159), .A3(n158), .ZN(n169) );
  nd02d1 U324 ( .A1(n162), .A2(n161), .ZN(n168) );
  inv0d1 U325 ( .I(N161), .ZN(n163) );
  inv0d1 U326 ( .I(n347), .ZN(n182) );
  nd02d1 U327 ( .A1(n129), .A2(n53), .ZN(n164) );
  nd03d0 U328 ( .A1(n166), .A2(n165), .A3(n164), .ZN(n167) );
  an02d1 U329 ( .A1(N117), .A2(n224), .Z(n175) );
  nr02d0 U330 ( .A1(n175), .A2(n174), .ZN(n191) );
  an02d1 U331 ( .A1(n177), .A2(n176), .Z(n190) );
  inv0d1 U332 ( .I(n178), .ZN(n184) );
  an02d1 U333 ( .A1(N165), .A2(n182), .Z(n183) );
  nr04d0 U334 ( .A1(n185), .A2(n184), .A3(n6), .A4(n183), .ZN(n186) );
  an02d1 U335 ( .A1(N116), .A2(n224), .Z(n194) );
  nr02d0 U336 ( .A1(n194), .A2(n193), .ZN(n211) );
  an02d1 U337 ( .A1(n196), .A2(n195), .Z(n210) );
  nd02d1 U338 ( .A1(n198), .A2(n197), .ZN(n205) );
  nd02d1 U339 ( .A1(n105), .A2(n53), .ZN(n199) );
  nd03d0 U340 ( .A1(n201), .A2(n200), .A3(n199), .ZN(n202) );
  nr02d0 U341 ( .A1(n205), .A2(n202), .ZN(n207) );
  nd02d1 U342 ( .A1(n13), .A2(n14), .ZN(n237) );
  an02d1 U343 ( .A1(N118), .A2(n224), .Z(n214) );
  nr02d0 U344 ( .A1(n214), .A2(n213), .ZN(n223) );
  an02d1 U345 ( .A1(n216), .A2(n215), .Z(n222) );
  nd02d1 U346 ( .A1(n218), .A2(n217), .ZN(n220) );
  nr03d0 U347 ( .A1(n220), .A2(n219), .A3(n52), .ZN(n221) );
  nd03d0 U348 ( .A1(n223), .A2(n222), .A3(n221), .ZN(n375) );
  an02d1 U349 ( .A1(N119), .A2(n224), .Z(n227) );
  nr02d0 U350 ( .A1(n227), .A2(n226), .ZN(n236) );
  an02d1 U351 ( .A1(n229), .A2(n228), .Z(n235) );
  nd02d1 U352 ( .A1(n231), .A2(n230), .ZN(n233) );
  nr03d0 U353 ( .A1(n233), .A2(n232), .A3(n51), .ZN(n234) );
  nd03d0 U354 ( .A1(n236), .A2(n235), .A3(n234), .ZN(n376) );
  nr03d0 U355 ( .A1(n237), .A2(n375), .A3(n376), .ZN(n360) );
  nr02d0 U356 ( .A1(n238), .A2(n53), .ZN(n241) );
  nr02d0 U357 ( .A1(n348), .A2(n239), .ZN(n240) );
  nr02d0 U358 ( .A1(n243), .A2(n242), .ZN(n249) );
  nr02d0 U359 ( .A1(n252), .A2(n53), .ZN(n255) );
  nr02d0 U360 ( .A1(n348), .A2(n253), .ZN(n254) );
  nr02d0 U361 ( .A1(n257), .A2(n256), .ZN(n265) );
  nr02d0 U362 ( .A1(n258), .A2(n338), .ZN(n263) );
  nr02d0 U363 ( .A1(n259), .A2(n347), .ZN(n261) );
  nr02d0 U364 ( .A1(n38), .A2(Oprnd_B[13]), .ZN(n260) );
  nr04d0 U365 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(n264) );
  an04d1 U366 ( .A1(n267), .A2(n266), .A3(n265), .A4(n264), .Z(n371) );
  nr02d0 U367 ( .A1(n268), .A2(n53), .ZN(n271) );
  nr02d0 U368 ( .A1(n348), .A2(n269), .ZN(n270) );
  nr02d0 U369 ( .A1(n273), .A2(n272), .ZN(n281) );
  nr02d0 U370 ( .A1(n274), .A2(n338), .ZN(n279) );
  nr02d0 U371 ( .A1(n275), .A2(n347), .ZN(n277) );
  nr02d0 U372 ( .A1(n38), .A2(Oprnd_B[12]), .ZN(n276) );
  nr04d0 U373 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .ZN(n280) );
  an04d1 U374 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .Z(n370) );
  an02d1 U375 ( .A1(n285), .A2(n284), .Z(n298) );
  nd02d1 U376 ( .A1(n287), .A2(n286), .ZN(n296) );
  mx02d0 U377 ( .I0(n74), .I1(n54), .S(Oprnd_B[11]), .Z(n288) );
  nr02d0 U378 ( .A1(n288), .A2(n53), .ZN(n291) );
  nr02d0 U379 ( .A1(n289), .A2(n348), .ZN(n290) );
  nd02d1 U380 ( .A1(n294), .A2(n293), .ZN(n295) );
  nr02d0 U381 ( .A1(n296), .A2(n295), .ZN(n297) );
  an02d1 U382 ( .A1(n370), .A2(n15), .Z(n358) );
  nd02d1 U383 ( .A1(n302), .A2(n301), .ZN(n305) );
  nr02d0 U384 ( .A1(n305), .A2(n304), .ZN(n312) );
  nr02d0 U385 ( .A1(n307), .A2(n306), .ZN(n308) );
  an03d1 U386 ( .A1(n310), .A2(n309), .A3(n308), .Z(n311) );
  nd02d1 U387 ( .A1(n312), .A2(n311), .ZN(n364) );
  nd02d1 U388 ( .A1(n314), .A2(n313), .ZN(n317) );
  nr02d0 U389 ( .A1(n317), .A2(n316), .ZN(n324) );
  nr02d0 U390 ( .A1(n319), .A2(n318), .ZN(n320) );
  an03d1 U391 ( .A1(n322), .A2(n321), .A3(n320), .Z(n323) );
  nd02d1 U392 ( .A1(n326), .A2(n325), .ZN(n329) );
  nr02d0 U393 ( .A1(n329), .A2(n328), .ZN(n336) );
  nr02d0 U394 ( .A1(n331), .A2(n330), .ZN(n332) );
  an03d1 U395 ( .A1(n334), .A2(n333), .A3(n332), .Z(n335) );
  nd02d1 U396 ( .A1(n336), .A2(n335), .ZN(n366) );
  nd02d1 U397 ( .A1(n340), .A2(n339), .ZN(n345) );
  nr02d0 U398 ( .A1(n345), .A2(n344), .ZN(n355) );
  nr02d0 U399 ( .A1(n350), .A2(n349), .ZN(n351) );
  an03d1 U400 ( .A1(n353), .A2(n352), .A3(n351), .Z(n354) );
  nd02d1 U401 ( .A1(n355), .A2(n354), .ZN(n368) );
  nr03d0 U402 ( .A1(n356), .A2(n366), .A3(n368), .ZN(n357) );
  nr02d0 U403 ( .A1(n36), .A2(n57), .ZN(Result[7]) );
  nr02d0 U404 ( .A1(n365), .A2(n57), .ZN(Result[8]) );
  nr02d0 U405 ( .A1(n367), .A2(n57), .ZN(Result[9]) );
  nr02d0 U406 ( .A1(n369), .A2(n57), .ZN(Result[10]) );
  nr02d0 U407 ( .A1(n15), .A2(n57), .ZN(Result[11]) );
  nr02d0 U408 ( .A1(n370), .A2(n57), .ZN(Result[12]) );
  nr02d0 U409 ( .A1(n371), .A2(n57), .ZN(Result[13]) );
  nr02d0 U410 ( .A1(n372), .A2(n57), .ZN(Result[14]) );
  inv0d1 U411 ( .I(ALU_OP[1]), .ZN(n394) );
  inv0d1 U412 ( .I(n373), .ZN(n377) );
  inv0d1 U413 ( .I(n374), .ZN(n378) );
endmodule


module PCI_FIFO_1 ( fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, 
        fifo_push_req_n, fifo_pop_req_n, fifo_data_in, push_empty_fifo, 
        push_ae_fifo, push_hf_fifo, push_af_fifo, push_full_fifo, 
        push_error_fifo, pop_empty_fifo, pop_ae_fifo, pop_hf_fifo, pop_af_fifo, 
        pop_full_fifo, pop_error_fifo, data_out_fifo, test_si1, test_si2, 
        test_se, test_so1, test_so2 );
  input [31:0] fifo_data_in;
  output [31:0] data_out_fifo;
  input fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, fifo_push_req_n,
         fifo_pop_req_n, test_si1, test_si2, test_se;
  output push_empty_fifo, push_ae_fifo, push_hf_fifo, push_af_fifo,
         push_full_fifo, push_error_fifo, pop_empty_fifo, pop_ae_fifo,
         pop_hf_fifo, pop_af_fifo, pop_full_fifo, pop_error_fifo, test_so1,
         test_so2;
  wire   we_n, wr_addr_5_, wr_addr_4_, wr_addr_3_, wr_addr_2_, wr_addr_1_,
         wr_addr_0_, rd_addr_5_, rd_addr_4_, rd_addr_3_, rd_addr_2_,
         rd_addr_1_, rd_addr_0_, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92;

  ram8x64 PCI_FIFO_RAM_1 ( .A1({wr_addr_5_, wr_addr_4_, wr_addr_3_, wr_addr_2_, 
        wr_addr_1_, wr_addr_0_}), .A2({rd_addr_5_, rd_addr_4_, rd_addr_3_, 
        rd_addr_2_, rd_addr_1_, rd_addr_0_}), .I1(fifo_data_in[7:0]), .O1({
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[7:0]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram8x64 PCI_FIFO_RAM_2 ( .A1({wr_addr_5_, wr_addr_4_, wr_addr_3_, wr_addr_2_, 
        wr_addr_1_, wr_addr_0_}), .A2({rd_addr_5_, rd_addr_4_, rd_addr_3_, 
        rd_addr_2_, rd_addr_1_, rd_addr_0_}), .I1(fifo_data_in[15:8]), .O1({
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[15:8]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram8x64 PCI_FIFO_RAM_3 ( .A1({wr_addr_5_, wr_addr_4_, wr_addr_3_, wr_addr_2_, 
        wr_addr_1_, wr_addr_0_}), .A2({rd_addr_5_, rd_addr_4_, rd_addr_3_, 
        rd_addr_2_, rd_addr_1_, rd_addr_0_}), .I1(fifo_data_in[23:16]), .O1({
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[23:16]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram8x64 PCI_FIFO_RAM_4 ( .A1({wr_addr_5_, wr_addr_4_, wr_addr_3_, wr_addr_2_, 
        wr_addr_1_, wr_addr_0_}), .A2({rd_addr_5_, rd_addr_4_, rd_addr_3_, 
        rd_addr_2_, rd_addr_1_, rd_addr_0_}), .I1(fifo_data_in[31:24]), .O1({
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[31:24]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  PCI_FIFO_1_DW_fifoctl_s2_sf_0 PCI_FIFO_CTL ( .clk_push(fifo_clk_push), 
        .clk_pop(fifo_clk_pop), .rst_n(fifo_rst_n), .push_req_n(
        fifo_push_req_n), .pop_req_n(fifo_pop_req_n), .we_n(we_n), 
        .push_empty(push_empty_fifo), .push_ae(push_ae_fifo), .push_hf(
        push_hf_fifo), .push_af(push_af_fifo), .push_full(push_full_fifo), 
        .push_error(push_error_fifo), .pop_empty(pop_empty_fifo), .pop_ae(
        pop_ae_fifo), .pop_hf(pop_hf_fifo), .pop_af(pop_af_fifo), .pop_full(
        pop_full_fifo), .pop_error(pop_error_fifo), .wr_addr({wr_addr_5_, 
        wr_addr_4_, wr_addr_3_, wr_addr_2_, wr_addr_1_, wr_addr_0_}), 
        .rd_addr({rd_addr_5_, rd_addr_4_, rd_addr_3_, rd_addr_2_, rd_addr_1_, 
        rd_addr_0_}), .push_word_count({SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85}), .pop_word_count({
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92}), .test(test_mode), .test_si1(test_si1), 
        .test_si2(test_si2), .test_se(test_se), .test_so2(test_so2), 
        .test_so1(test_so1) );
endmodule


module PCI_FIFO_0 ( fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, 
        fifo_push_req_n, fifo_pop_req_n, fifo_data_in, push_empty_fifo, 
        push_ae_fifo, push_hf_fifo, push_af_fifo, push_full_fifo, 
        push_error_fifo, pop_empty_fifo, pop_ae_fifo, pop_hf_fifo, pop_af_fifo, 
        pop_full_fifo, pop_error_fifo, data_out_fifo, test_si1, test_si2, 
        test_se, test_so1, test_so2 );
  input [31:0] fifo_data_in;
  output [31:0] data_out_fifo;
  input fifo_clk_push, fifo_clk_pop, fifo_rst_n, test_mode, fifo_push_req_n,
         fifo_pop_req_n, test_si1, test_si2, test_se;
  output push_empty_fifo, push_ae_fifo, push_hf_fifo, push_af_fifo,
         push_full_fifo, push_error_fifo, pop_empty_fifo, pop_ae_fifo,
         pop_hf_fifo, pop_af_fifo, pop_full_fifo, pop_error_fifo, test_so1,
         test_so2;
  wire   we_n, SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92;
  wire   [5:0] wr_addr;
  wire   [5:0] rd_addr;

  ram8x64 PCI_FIFO_RAM_1 ( .A1(wr_addr), .A2(rd_addr), .I1(fifo_data_in[7:0]), 
        .O1({SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[7:0]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram8x64 PCI_FIFO_RAM_2 ( .A1(wr_addr), .A2(rd_addr), .I1(fifo_data_in[15:8]), 
        .O1({SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[15:8]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram8x64 PCI_FIFO_RAM_3 ( .A1(wr_addr), .A2(rd_addr), .I1(fifo_data_in[23:16]), .O1({SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[23:16]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  ram8x64 PCI_FIFO_RAM_4 ( .A1(wr_addr), .A2(rd_addr), .I1(fifo_data_in[31:24]), .O1({SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78}), .I2({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .O2(data_out_fifo[31:24]), .CE1(
        fifo_clk_push), .CE2(fifo_clk_pop), .OEB1(1'b1), .OEB2(1'b0), .CSB1(
        1'b0), .CSB2(1'b0), .WEB1(we_n), .WEB2(1'b1) );
  PCI_FIFO_0_DW_fifoctl_s2_sf_0 PCI_FIFO_CTL ( .clk_push(fifo_clk_push), 
        .clk_pop(fifo_clk_pop), .rst_n(fifo_rst_n), .push_req_n(
        fifo_push_req_n), .pop_req_n(fifo_pop_req_n), .we_n(we_n), 
        .push_empty(push_empty_fifo), .push_ae(push_ae_fifo), .push_hf(
        push_hf_fifo), .push_af(push_af_fifo), .push_full(push_full_fifo), 
        .push_error(push_error_fifo), .pop_empty(pop_empty_fifo), .pop_ae(
        pop_ae_fifo), .pop_hf(pop_hf_fifo), .pop_af(pop_af_fifo), .pop_full(
        pop_full_fifo), .pop_error(pop_error_fifo), .wr_addr(wr_addr), 
        .rd_addr(rd_addr), .push_word_count({SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85}), .pop_word_count({
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92}), .test(test_mode), .test_si1(test_si1), 
        .test_si2(test_si2), .test_se(test_se), .test_so2(test_so2), 
        .test_so1(test_so1) );
endmodule


module PCI_CORE ( pclk, pci_rst_n, pidsel, pgnt_n, pad_in, pad_out, pad_en, 
        ppar_in, ppar_out, ppar_en, pc_be_in, pc_be_out, pc_be_en, pframe_n_in, 
        pframe_n_out, pframe_n_en, ptrdy_n_in, ptrdy_n_out, ptrdy_n_en, 
        pirdy_n_in, pirdy_n_out, pirdy_n_en, pdevsel_n_in, pdevsel_n_out, 
        pdevsel_n_en, pstop_n_in, pstop_n_out, pstop_n_en, pperr_n_in, 
        pperr_n_out, pperr_n_en, pserr_n_in, pserr_n_out, pserr_n_en, preq_n, 
        pm66en, read_data, write_data, read_push, read_full, write_pop, 
        write_empty, cmd_valid, cmd, cmd_in_valid, cmd_in, test_se, test_si1, 
        test_si2 );
  input [15:0] pad_in;
  output [15:0] pad_out;
  input [3:0] pc_be_in;
  output [3:0] pc_be_out;
  output [31:0] read_data;
  input [31:0] write_data;
  output [3:0] cmd;
  input [3:0] cmd_in;
  input pclk, pci_rst_n, pidsel, pgnt_n, ppar_in, pframe_n_in, ptrdy_n_in,
         pirdy_n_in, pdevsel_n_in, pstop_n_in, pperr_n_in, pserr_n_in, pm66en,
         read_full, write_empty, cmd_in_valid, test_se, test_si1, test_si2;
  output pad_en, ppar_out, ppar_en, pc_be_en, pframe_n_out, pframe_n_en,
         ptrdy_n_out, ptrdy_n_en, pirdy_n_out, pirdy_n_en, pdevsel_n_out,
         pdevsel_n_en, pstop_n_out, pstop_n_en, pperr_n_out, pperr_n_en,
         pserr_n_out, pserr_n_en, preq_n, read_push, write_pop, cmd_valid;
  wire   N45, N46, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N118, N119,
         N120, N121, N122, N123, N124, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n1, n214;
  wire   [79:0] mega_shift;

  sdcrn1 d_out_p_bus_reg_3_ ( .D(N75), .SD(ppar_en), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .QN(N46) );
  sdcrn1 d_out_p_bus_reg_0_ ( .D(N72), .SD(cmd[3]), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .QN(N45) );
  an02d1 U143 ( .A1(n214), .A2(n139), .Z(N73) );
  an03d1 U150 ( .A1(read_full), .A2(cmd_in[0]), .A3(n172), .Z(n170) );
  an02d1 U160 ( .A1(n189), .A2(n190), .Z(n181) );
  an02d1 U161 ( .A1(n191), .A2(n175), .Z(n178) );
  an04d1 U165 ( .A1(n197), .A2(n198), .A3(n199), .A4(n200), .Z(n191) );
  an04d1 U168 ( .A1(n198), .A2(n203), .A3(pirdy_n_in), .A4(n195), .Z(n202) );
  an03d1 U172 ( .A1(n203), .A2(n206), .A3(n196), .Z(n211) );
  an03d1 U173 ( .A1(pirdy_n_in), .A2(n207), .A3(n212), .Z(n196) );
  an04d1 U174 ( .A1(n206), .A2(n207), .A3(n195), .A4(n213), .Z(n208) );
  aor22d1 U183 ( .A1(pad_in[1]), .A2(n130), .B1(pad_in[9]), .B2(n131), .Z(
        read_data[9]) );
  aor22d1 U184 ( .A1(pad_in[0]), .A2(n130), .B1(pad_in[8]), .B2(n131), .Z(
        read_data[8]) );
  an12d1 U185 ( .A2(pad_in[7]), .A1(n132), .Z(read_data[7]) );
  an12d1 U186 ( .A2(pad_in[6]), .A1(n132), .Z(read_data[6]) );
  an12d1 U187 ( .A2(pad_in[5]), .A1(n132), .Z(read_data[5]) );
  an12d1 U188 ( .A2(pad_in[4]), .A1(n132), .Z(read_data[4]) );
  an12d1 U189 ( .A2(pad_in[3]), .A1(n132), .Z(read_data[3]) );
  an12d1 U190 ( .A2(pad_in[15]), .A1(n133), .Z(read_data[31]) );
  an12d1 U191 ( .A2(pad_in[14]), .A1(n133), .Z(read_data[30]) );
  an12d1 U192 ( .A2(pad_in[2]), .A1(n132), .Z(read_data[2]) );
  an12d1 U193 ( .A2(pad_in[13]), .A1(n133), .Z(read_data[29]) );
  an12d1 U194 ( .A2(pad_in[12]), .A1(n133), .Z(read_data[28]) );
  an12d1 U195 ( .A2(pad_in[11]), .A1(n133), .Z(read_data[27]) );
  an12d1 U196 ( .A2(pad_in[10]), .A1(n133), .Z(read_data[26]) );
  an12d1 U197 ( .A2(pad_in[9]), .A1(n133), .Z(read_data[25]) );
  an12d1 U198 ( .A2(pad_in[8]), .A1(n133), .Z(read_data[24]) );
  nr02d0 U199 ( .A1(n134), .A2(n130), .ZN(n133) );
  aor22d1 U200 ( .A1(n134), .A2(pad_in[7]), .B1(n135), .B2(pad_in[15]), .Z(
        read_data[23]) );
  aor22d1 U201 ( .A1(n134), .A2(pad_in[6]), .B1(n135), .B2(pad_in[14]), .Z(
        read_data[22]) );
  aor22d1 U202 ( .A1(n134), .A2(pad_in[5]), .B1(n135), .B2(pad_in[13]), .Z(
        read_data[21]) );
  aor22d1 U203 ( .A1(n134), .A2(pad_in[4]), .B1(n135), .B2(pad_in[12]), .Z(
        read_data[20]) );
  an12d1 U204 ( .A2(pad_in[1]), .A1(n132), .Z(read_data[1]) );
  aor22d1 U205 ( .A1(n134), .A2(pad_in[3]), .B1(n135), .B2(pad_in[11]), .Z(
        read_data[19]) );
  aor22d1 U206 ( .A1(n134), .A2(pad_in[2]), .B1(n135), .B2(pad_in[10]), .Z(
        read_data[18]) );
  aor22d1 U207 ( .A1(n134), .A2(pad_in[1]), .B1(n135), .B2(pad_in[9]), .Z(
        read_data[17]) );
  aor22d1 U208 ( .A1(n134), .A2(pad_in[0]), .B1(n135), .B2(pad_in[8]), .Z(
        read_data[16]) );
  aor22d1 U209 ( .A1(pad_in[7]), .A2(n130), .B1(pad_in[15]), .B2(n131), .Z(
        read_data[15]) );
  aor22d1 U210 ( .A1(pad_in[6]), .A2(n130), .B1(pad_in[14]), .B2(n131), .Z(
        read_data[14]) );
  aor22d1 U211 ( .A1(pad_in[5]), .A2(n130), .B1(pad_in[13]), .B2(n131), .Z(
        read_data[13]) );
  aor22d1 U212 ( .A1(pad_in[4]), .A2(n130), .B1(pad_in[12]), .B2(n131), .Z(
        read_data[12]) );
  aor22d1 U213 ( .A1(pad_in[3]), .A2(n130), .B1(pad_in[11]), .B2(n131), .Z(
        read_data[11]) );
  aor22d1 U214 ( .A1(pad_in[2]), .A2(n130), .B1(pad_in[10]), .B2(n131), .Z(
        read_data[10]) );
  an12d1 U216 ( .A2(pad_in[0]), .A1(n132), .Z(read_data[0]) );
  nr02d0 U217 ( .A1(n131), .A2(n135), .ZN(n132) );
  aor21d1 U219 ( .B1(write_data[18]), .B2(n139), .A(n140), .Z(N94) );
  aor21d1 U220 ( .B1(write_data[17]), .B2(n139), .A(n141), .Z(N93) );
  aor21d1 U221 ( .B1(write_data[16]), .B2(n139), .A(n140), .Z(N92) );
  aor211d1 U222 ( .C1(write_data[15]), .C2(n139), .A(n142), .B(n143), .Z(N91)
         );
  aor21d1 U223 ( .B1(write_data[13]), .B2(n139), .A(n141), .Z(N89) );
  nd04d0 U224 ( .A1(n146), .A2(n147), .A3(n148), .A4(n144), .ZN(N88) );
  aor21d1 U225 ( .B1(write_data[11]), .B2(n139), .A(n141), .Z(N87) );
  aor211d1 U226 ( .C1(write_data[10]), .C2(n139), .A(n149), .B(n150), .Z(N86)
         );
  aor21d1 U227 ( .B1(write_data[9]), .B2(n139), .A(n141), .Z(N85) );
  aor21d1 U228 ( .B1(write_data[8]), .B2(n139), .A(n150), .Z(N84) );
  aor21d1 U229 ( .B1(write_data[7]), .B2(n139), .A(n141), .Z(N83) );
  nd04d0 U230 ( .A1(n151), .A2(n152), .A3(n153), .A4(n148), .ZN(N82) );
  nr03d0 U231 ( .A1(n142), .A2(n140), .A3(n143), .ZN(n151) );
  nr03d0 U232 ( .A1(n154), .A2(n155), .A3(n156), .ZN(n142) );
  aor21d1 U233 ( .B1(write_data[5]), .B2(n139), .A(n141), .Z(N81) );
  aor211d1 U234 ( .C1(write_data[4]), .C2(n139), .A(n140), .B(n157), .Z(N80)
         );
  aor21d1 U235 ( .B1(write_data[3]), .B2(n139), .A(n141), .Z(N79) );
  aor211d1 U236 ( .C1(write_data[2]), .C2(n139), .A(n143), .B(n158), .Z(N78)
         );
  nd03d0 U237 ( .A1(n148), .A2(n144), .A3(n159), .ZN(n158) );
  nr03d0 U238 ( .A1(n155), .A2(write_empty), .A3(n156), .ZN(n149) );
  aor21d1 U239 ( .B1(write_data[1]), .B2(n139), .A(n141), .Z(N77) );
  nd04d0 U240 ( .A1(n160), .A2(n159), .A3(n144), .A4(n161), .ZN(N76) );
  aor21d1 U241 ( .B1(n139), .B2(cmd_in[3]), .A(n141), .Z(N75) );
  nd04d0 U243 ( .A1(n164), .A2(n163), .A3(n162), .A4(n165), .ZN(n144) );
  nd03d0 U245 ( .A1(read_full), .A2(n167), .A3(n168), .ZN(n161) );
  nr03d0 U246 ( .A1(n154), .A2(n155), .A3(n169), .ZN(n168) );
  nd04d0 U247 ( .A1(n171), .A2(n145), .A3(n159), .A4(n147), .ZN(n157) );
  nr04d0 U248 ( .A1(n154), .A2(n169), .A3(n155), .A4(read_full), .ZN(n164) );
  nd03d0 U249 ( .A1(n169), .A2(n165), .A3(n170), .ZN(n159) );
  nd03d0 U250 ( .A1(cmd_in_valid), .A2(cmd_in[3]), .A3(n170), .ZN(n145) );
  nr03d0 U251 ( .A1(n214), .A2(write_empty), .A3(cmd_in[2]), .ZN(n172) );
  nr03d0 U252 ( .A1(n214), .A2(write_empty), .A3(n156), .ZN(n143) );
  nd03d0 U253 ( .A1(n167), .A2(n169), .A3(read_full), .ZN(n156) );
  nr03d0 U254 ( .A1(n162), .A2(n163), .A3(n165), .ZN(n167) );
  aor22d1 U255 ( .A1(write_data[31]), .A2(n1), .B1(write_data[15]), .B2(n155), 
        .Z(N141) );
  aor22d1 U256 ( .A1(write_data[30]), .A2(n1), .B1(write_data[14]), .B2(n155), 
        .Z(N140) );
  aor22d1 U257 ( .A1(write_data[29]), .A2(n1), .B1(write_data[13]), .B2(n155), 
        .Z(N139) );
  aor22d1 U258 ( .A1(write_data[28]), .A2(n1), .B1(write_data[12]), .B2(n155), 
        .Z(N138) );
  aor22d1 U259 ( .A1(write_data[27]), .A2(n1), .B1(write_data[11]), .B2(n155), 
        .Z(N137) );
  aor22d1 U260 ( .A1(write_data[26]), .A2(n1), .B1(write_data[10]), .B2(n155), 
        .Z(N136) );
  aor22d1 U261 ( .A1(write_data[25]), .A2(n214), .B1(write_data[9]), .B2(n155), 
        .Z(N135) );
  aor22d1 U262 ( .A1(write_data[24]), .A2(n214), .B1(write_data[8]), .B2(n155), 
        .Z(N134) );
  aor22d1 U263 ( .A1(write_data[23]), .A2(n214), .B1(write_data[7]), .B2(n155), 
        .Z(N133) );
  aor22d1 U264 ( .A1(write_data[22]), .A2(n214), .B1(write_data[6]), .B2(n155), 
        .Z(N132) );
  aor22d1 U265 ( .A1(write_data[21]), .A2(n214), .B1(write_data[5]), .B2(n155), 
        .Z(N131) );
  aor22d1 U266 ( .A1(write_data[20]), .A2(n1), .B1(write_data[4]), .B2(n155), 
        .Z(N130) );
  aor22d1 U267 ( .A1(write_data[19]), .A2(n214), .B1(write_data[3]), .B2(n155), 
        .Z(N129) );
  aor22d1 U268 ( .A1(write_data[18]), .A2(n214), .B1(write_data[2]), .B2(n155), 
        .Z(N128) );
  aor22d1 U269 ( .A1(write_data[17]), .A2(n1), .B1(write_data[1]), .B2(n155), 
        .Z(N127) );
  aor22d1 U270 ( .A1(write_data[16]), .A2(n214), .B1(write_data[0]), .B2(n155), 
        .Z(N126) );
  aor221d1 U271 ( .B1(pad_in[6]), .B2(n173), .C1(n174), .C2(n175), .A(n176), 
        .Z(N124) );
  aor221d1 U272 ( .B1(n175), .B2(n177), .C1(pad_in[5]), .C2(n173), .A(n178), 
        .Z(N123) );
  aor221d1 U273 ( .B1(n175), .B2(n179), .C1(pad_in[4]), .C2(n173), .A(n180), 
        .Z(N122) );
  aor221d1 U274 ( .B1(n175), .B2(n177), .C1(pad_in[3]), .C2(n173), .A(n180), 
        .Z(N121) );
  aor221d1 U275 ( .B1(n175), .B2(n185), .C1(pad_in[2]), .C2(n173), .A(n180), 
        .Z(N120) );
  nr02d0 U276 ( .A1(n186), .A2(n187), .ZN(n180) );
  aor221d1 U277 ( .B1(n175), .B2(n188), .C1(pad_in[1]), .C2(n173), .A(n178), 
        .Z(N119) );
  aor21d1 U278 ( .B1(pad_in[0]), .B2(n173), .A(n176), .Z(N118) );
  aor21d1 U279 ( .B1(n175), .B2(n185), .A(n178), .Z(n176) );
  aor31d1 U280 ( .B1(n192), .B2(n186), .B3(n193), .A(n187), .Z(n173) );
  nr03d0 U281 ( .A1(n194), .A2(n191), .A3(n174), .ZN(n193) );
  nd04d0 U282 ( .A1(pframe_n_in), .A2(pdevsel_n_in), .A3(n195), .A4(n196), 
        .ZN(n189) );
  nr04d0 U283 ( .A1(pidsel), .A2(pgnt_n), .A3(pframe_n_in), .A4(pdevsel_n_in), 
        .ZN(n200) );
  nr03d0 U284 ( .A1(pperr_n_in), .A2(ptrdy_n_in), .A3(pserr_n_in), .ZN(n199)
         );
  nr04d0 U285 ( .A1(n204), .A2(n205), .A3(n206), .A4(n207), .ZN(n201) );
  nd03d0 U286 ( .A1(n208), .A2(n197), .A3(pdevsel_n_in), .ZN(n186) );
  nd03d0 U287 ( .A1(n183), .A2(n182), .A3(n190), .ZN(n185) );
  nd03d0 U288 ( .A1(n209), .A2(n210), .A3(n211), .ZN(n190) );
  nr03d0 U289 ( .A1(pm66en), .A2(ptrdy_n_in), .A3(pperr_n_in), .ZN(n212) );
  nd03d0 U290 ( .A1(pirdy_n_in), .A2(n203), .A3(n208), .ZN(n183) );
  nr03d0 U291 ( .A1(n205), .A2(n198), .A3(n204), .ZN(n213) );
  nr02d0 U292 ( .A1(n210), .A2(n209), .ZN(n195) );
  PCI_CORE_DW_mult_uns_0 mult_43_L43980_C240_I4 ( .a(mega_shift[15:8]), .b(
        mega_shift[7:0]), .product({N205, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190}) );
  PCI_CORE_DW_mult_uns_1 mult_43_L43980_C240_I3 ( .a(mega_shift[31:24]), .b(
        mega_shift[23:16]), .product({N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174}) );
  PCI_CORE_DW_mult_uns_2 mult_43_L43980_C240_I2 ( .a(mega_shift[47:40]), .b(
        mega_shift[39:32]), .product({N173, N172, N171, N170, N169, N168, N167, 
        N166, N165, N164, N163, N162, N161, N160, N159, N158}) );
  PCI_CORE_DW_mult_uns_3 mult_43_L43980_C240 ( .a(mega_shift[63:56]), .b(
        mega_shift[55:48]), .product({N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142}) );
  sdcrq1 d_out_i_bus_reg_1_ ( .D(N119), .SD(read_push), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(write_pop) );
  sdcrq1 d_out_i_bus_reg_0_ ( .D(N118), .SD(test_si1), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(read_push) );
  sdcrq1 mega_shift_reg_1__15_ ( .D(N173), .SD(mega_shift[62]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[63]) );
  sdcrq1 mega_shift_reg_1__14_ ( .D(N172), .SD(mega_shift[61]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[62]) );
  sdcrq1 mega_shift_reg_1__13_ ( .D(N171), .SD(mega_shift[60]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[61]) );
  sdcrq1 mega_shift_reg_1__12_ ( .D(N170), .SD(mega_shift[59]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[60]) );
  sdcrq1 mega_shift_reg_1__11_ ( .D(N169), .SD(mega_shift[58]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[59]) );
  sdcrq1 mega_shift_reg_1__10_ ( .D(N168), .SD(mega_shift[57]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[58]) );
  sdcrq1 mega_shift_reg_1__9_ ( .D(N167), .SD(mega_shift[56]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[57]) );
  sdcrq1 mega_shift_reg_1__8_ ( .D(N166), .SD(mega_shift[55]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[56]) );
  sdcrq1 mega_shift_reg_1__7_ ( .D(N165), .SD(mega_shift[54]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[55]) );
  sdcrq1 mega_shift_reg_1__6_ ( .D(N164), .SD(mega_shift[53]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[54]) );
  sdcrq1 mega_shift_reg_1__5_ ( .D(N163), .SD(mega_shift[52]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[53]) );
  sdcrq1 mega_shift_reg_1__4_ ( .D(N162), .SD(mega_shift[51]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[52]) );
  sdcrq1 mega_shift_reg_1__3_ ( .D(N161), .SD(mega_shift[50]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[51]) );
  sdcrq1 mega_shift_reg_1__2_ ( .D(N160), .SD(mega_shift[49]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[50]) );
  sdcrq1 mega_shift_reg_1__1_ ( .D(N159), .SD(mega_shift[48]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[49]) );
  sdcrq1 mega_shift_reg_1__0_ ( .D(N158), .SD(mega_shift[79]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[48]) );
  sdcrq1 mega_shift_reg_2__15_ ( .D(N189), .SD(mega_shift[46]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[47]) );
  sdcrq1 mega_shift_reg_2__14_ ( .D(N188), .SD(mega_shift[45]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[46]) );
  sdcrq1 mega_shift_reg_2__13_ ( .D(N187), .SD(mega_shift[44]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[45]) );
  sdcrq1 mega_shift_reg_2__12_ ( .D(N186), .SD(mega_shift[43]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[44]) );
  sdcrq1 mega_shift_reg_2__11_ ( .D(N185), .SD(mega_shift[42]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[43]) );
  sdcrq1 mega_shift_reg_2__10_ ( .D(N184), .SD(mega_shift[41]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[42]) );
  sdcrq1 mega_shift_reg_2__9_ ( .D(N183), .SD(mega_shift[40]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[41]) );
  sdcrq1 mega_shift_reg_2__8_ ( .D(N182), .SD(mega_shift[39]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[40]) );
  sdcrq1 mega_shift_reg_2__7_ ( .D(N181), .SD(mega_shift[38]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[39]) );
  sdcrq1 mega_shift_reg_2__6_ ( .D(N180), .SD(mega_shift[37]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[38]) );
  sdcrq1 mega_shift_reg_2__5_ ( .D(N179), .SD(mega_shift[36]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[37]) );
  sdcrq1 mega_shift_reg_2__4_ ( .D(N178), .SD(mega_shift[35]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[36]) );
  sdcrq1 mega_shift_reg_2__3_ ( .D(N177), .SD(mega_shift[34]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[35]) );
  sdcrq1 mega_shift_reg_2__2_ ( .D(N176), .SD(mega_shift[33]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[34]) );
  sdcrq1 mega_shift_reg_2__1_ ( .D(N175), .SD(mega_shift[32]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[33]) );
  sdcrq1 mega_shift_reg_2__0_ ( .D(N174), .SD(mega_shift[63]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[32]) );
  sdcrq1 mega_shift_reg_3__15_ ( .D(N205), .SD(mega_shift[30]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[31]) );
  sdcrq1 mega_shift_reg_3__14_ ( .D(N204), .SD(mega_shift[29]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[30]) );
  sdcrq1 mega_shift_reg_3__13_ ( .D(N203), .SD(mega_shift[28]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[29]) );
  sdcrq1 mega_shift_reg_3__12_ ( .D(N202), .SD(mega_shift[27]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[28]) );
  sdcrq1 mega_shift_reg_3__11_ ( .D(N201), .SD(mega_shift[26]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[27]) );
  sdcrq1 mega_shift_reg_3__10_ ( .D(N200), .SD(mega_shift[25]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[26]) );
  sdcrq1 mega_shift_reg_3__9_ ( .D(N199), .SD(mega_shift[24]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[25]) );
  sdcrq1 mega_shift_reg_3__8_ ( .D(N198), .SD(mega_shift[23]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[24]) );
  sdcrq1 mega_shift_reg_3__7_ ( .D(N197), .SD(mega_shift[22]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[23]) );
  sdcrq1 mega_shift_reg_3__6_ ( .D(N196), .SD(mega_shift[21]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[22]) );
  sdcrq1 mega_shift_reg_3__5_ ( .D(N195), .SD(mega_shift[20]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[21]) );
  sdcrq1 mega_shift_reg_3__4_ ( .D(N194), .SD(mega_shift[19]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[20]) );
  sdcrq1 mega_shift_reg_3__3_ ( .D(N193), .SD(mega_shift[18]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[19]) );
  sdcrq1 mega_shift_reg_3__2_ ( .D(N192), .SD(mega_shift[17]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[18]) );
  sdcrq1 mega_shift_reg_3__1_ ( .D(N191), .SD(mega_shift[16]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[17]) );
  sdcrq1 mega_shift_reg_3__0_ ( .D(N190), .SD(mega_shift[47]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[16]) );
  sdcrq1 mega_shift_reg_4__15_ ( .D(N141), .SD(mega_shift[14]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[15]) );
  sdcrq1 mega_shift_reg_4__14_ ( .D(N140), .SD(mega_shift[13]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[14]) );
  sdcrq1 mega_shift_reg_4__13_ ( .D(N139), .SD(mega_shift[12]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[13]) );
  sdcrq1 mega_shift_reg_4__12_ ( .D(N138), .SD(mega_shift[11]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[12]) );
  sdcrq1 mega_shift_reg_4__11_ ( .D(N137), .SD(mega_shift[10]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[11]) );
  sdcrq1 mega_shift_reg_4__10_ ( .D(N136), .SD(mega_shift[9]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[10]) );
  sdcrq1 mega_shift_reg_4__9_ ( .D(N135), .SD(mega_shift[8]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[9]) );
  sdcrq1 mega_shift_reg_4__8_ ( .D(N134), .SD(mega_shift[7]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[8]) );
  sdcrq1 mega_shift_reg_4__7_ ( .D(N133), .SD(mega_shift[6]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[7]) );
  sdcrq1 mega_shift_reg_4__6_ ( .D(N132), .SD(mega_shift[5]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[6]) );
  sdcrq1 mega_shift_reg_4__5_ ( .D(N131), .SD(mega_shift[4]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[5]) );
  sdcrq1 mega_shift_reg_4__4_ ( .D(N130), .SD(mega_shift[3]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[4]) );
  sdcrq1 mega_shift_reg_4__3_ ( .D(N129), .SD(mega_shift[2]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[3]) );
  sdcrq1 mega_shift_reg_4__2_ ( .D(N128), .SD(mega_shift[1]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[2]) );
  sdcrq1 mega_shift_reg_4__1_ ( .D(N127), .SD(mega_shift[0]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[1]) );
  sdcrq1 mega_shift_reg_4__0_ ( .D(N126), .SD(mega_shift[31]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[0]) );
  sdcrq1 d_out_i_bus_reg_6_ ( .D(N124), .SD(cmd[2]), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(cmd[3]) );
  sdcrq1 d_out_i_bus_reg_5_ ( .D(N123), .SD(cmd[1]), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(cmd[2]) );
  sdcrq1 d_out_i_bus_reg_4_ ( .D(N122), .SD(cmd[0]), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(cmd[1]) );
  sdcrq1 d_out_i_bus_reg_3_ ( .D(N121), .SD(cmd_valid), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(cmd[0]) );
  sdcrq1 d_out_i_bus_reg_2_ ( .D(N120), .SD(write_pop), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(cmd_valid) );
  sdcrq1 mega_shift_reg_0__14_ ( .D(N156), .SD(mega_shift[77]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[78]) );
  sdcrq1 mega_shift_reg_0__2_ ( .D(N144), .SD(mega_shift[65]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[66]) );
  sdcrq1 mega_shift_reg_0__1_ ( .D(N143), .SD(mega_shift[64]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[65]) );
  sdcrq1 mega_shift_reg_0__0_ ( .D(N142), .SD(pc_be_out[3]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[64]) );
  sdcrq1 mega_shift_reg_0__15_ ( .D(N157), .SD(mega_shift[78]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[79]) );
  sdcrq1 mega_shift_reg_0__13_ ( .D(N155), .SD(mega_shift[76]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[77]) );
  sdcrq1 mega_shift_reg_0__4_ ( .D(N146), .SD(mega_shift[67]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[68]) );
  sdcrq1 mega_shift_reg_0__3_ ( .D(N145), .SD(mega_shift[66]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[67]) );
  sdcrq1 mega_shift_reg_0__12_ ( .D(N154), .SD(mega_shift[75]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[76]) );
  sdcrq1 mega_shift_reg_0__11_ ( .D(N153), .SD(mega_shift[74]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[75]) );
  sdcrq1 mega_shift_reg_0__7_ ( .D(N149), .SD(mega_shift[70]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[71]) );
  sdcrq1 mega_shift_reg_0__6_ ( .D(N148), .SD(mega_shift[69]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[70]) );
  sdcrq1 mega_shift_reg_0__5_ ( .D(N147), .SD(mega_shift[68]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[69]) );
  sdcrq1 mega_shift_reg_0__10_ ( .D(N152), .SD(mega_shift[73]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[74]) );
  sdcrq1 mega_shift_reg_0__9_ ( .D(N151), .SD(mega_shift[72]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[73]) );
  sdcrq1 mega_shift_reg_0__8_ ( .D(N150), .SD(mega_shift[71]), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(mega_shift[72]) );
  sdcrq4 pad_out_buf_reg_0_ ( .D(mega_shift[64]), .SD(pad_en), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[0]) );
  sdcrq4 pad_out_buf_reg_1_ ( .D(mega_shift[65]), .SD(pad_out[0]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[1]) );
  sdcrq4 pad_out_buf_reg_2_ ( .D(mega_shift[66]), .SD(pad_out[1]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[2]) );
  sdcrq4 pad_out_buf_reg_3_ ( .D(mega_shift[67]), .SD(test_si2), .SC(test_se), 
        .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[3]) );
  sdcrq4 pad_out_buf_reg_4_ ( .D(mega_shift[68]), .SD(pad_out[3]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[4]) );
  sdcrq4 pad_out_buf_reg_5_ ( .D(mega_shift[69]), .SD(pad_out[4]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[5]) );
  sdcrq4 pad_out_buf_reg_6_ ( .D(mega_shift[70]), .SD(pad_out[5]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[6]) );
  sdcrq4 pad_out_buf_reg_7_ ( .D(mega_shift[71]), .SD(pad_out[6]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[7]) );
  sdcrq4 pad_out_buf_reg_8_ ( .D(mega_shift[72]), .SD(pad_out[7]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[8]) );
  sdcrq4 pad_out_buf_reg_9_ ( .D(mega_shift[73]), .SD(pad_out[8]), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[9]) );
  sdcrq4 pad_out_buf_reg_10_ ( .D(mega_shift[74]), .SD(pad_out[9]), .SC(
        test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[10]) );
  sdcrq4 pad_out_buf_reg_11_ ( .D(mega_shift[75]), .SD(pad_out[10]), .SC(
        test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[11]) );
  sdcrq4 pad_out_buf_reg_12_ ( .D(mega_shift[76]), .SD(pad_out[11]), .SC(
        test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[12]) );
  sdcrq4 pad_out_buf_reg_13_ ( .D(mega_shift[77]), .SD(pad_out[12]), .SC(
        test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[13]) );
  sdcrq4 pad_out_buf_reg_14_ ( .D(mega_shift[78]), .SD(pad_out[13]), .SC(
        test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[14]) );
  sdcrq4 pad_out_buf_reg_15_ ( .D(mega_shift[79]), .SD(pad_out[14]), .SC(
        test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pad_out[15]) );
  sdcrq4 pad_en_reg ( .D(N45), .SD(mega_shift[15]), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(pad_en) );
  sdcrq4 d_out_p_bus_reg_1_ ( .D(N73), .SD(N45), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(ppar_out) );
  sdcrq4 d_out_p_bus_reg_2_ ( .D(N74), .SD(ppar_out), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(ppar_en) );
  sdcrq4 pc_be_en_reg ( .D(N46), .SD(pad_out[15]), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(pc_be_en) );
  sdcrq4 d_out_p_bus_reg_4_ ( .D(N76), .SD(N46), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(pframe_n_out) );
  sdcrq4 d_out_p_bus_reg_5_ ( .D(N77), .SD(pframe_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pframe_n_en) );
  sdcrq4 d_out_p_bus_reg_6_ ( .D(N78), .SD(pframe_n_en), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(ptrdy_n_out) );
  sdcrq4 d_out_p_bus_reg_7_ ( .D(N79), .SD(ptrdy_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(ptrdy_n_en) );
  sdcrq4 d_out_p_bus_reg_8_ ( .D(N80), .SD(ptrdy_n_en), .SC(test_se), .CP(pclk), .CDN(pci_rst_n), .Q(pirdy_n_out) );
  sdcrq4 d_out_p_bus_reg_9_ ( .D(N81), .SD(pirdy_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pirdy_n_en) );
  sdcrq4 d_out_p_bus_reg_10_ ( .D(N82), .SD(pirdy_n_en), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pdevsel_n_out) );
  sdcrq4 d_out_p_bus_reg_11_ ( .D(N83), .SD(pdevsel_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pdevsel_n_en) );
  sdcrq4 d_out_p_bus_reg_12_ ( .D(N84), .SD(pdevsel_n_en), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pstop_n_out) );
  sdcrq4 d_out_p_bus_reg_13_ ( .D(N85), .SD(pstop_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pstop_n_en) );
  sdcrq4 d_out_p_bus_reg_14_ ( .D(N86), .SD(pstop_n_en), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pperr_n_out) );
  sdcrq4 d_out_p_bus_reg_15_ ( .D(N87), .SD(pperr_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pperr_n_en) );
  sdcrq4 d_out_p_bus_reg_16_ ( .D(N88), .SD(pperr_n_en), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pserr_n_out) );
  sdcrq4 d_out_p_bus_reg_17_ ( .D(N89), .SD(pserr_n_out), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pserr_n_en) );
  sdcrq4 d_out_p_bus_reg_18_ ( .D(N90), .SD(pserr_n_en), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(preq_n) );
  sdcrq4 d_out_p_bus_reg_19_ ( .D(N91), .SD(preq_n), .SC(test_se), .CP(pclk), 
        .CDN(pci_rst_n), .Q(pc_be_out[0]) );
  sdcrq4 d_out_p_bus_reg_20_ ( .D(N92), .SD(pc_be_out[0]), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pc_be_out[1]) );
  sdcrq4 d_out_p_bus_reg_21_ ( .D(N93), .SD(pc_be_out[1]), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pc_be_out[2]) );
  sdcrq4 d_out_p_bus_reg_22_ ( .D(N94), .SD(pc_be_out[2]), .SC(test_se), .CP(
        pclk), .CDN(pci_rst_n), .Q(pc_be_out[3]) );
  nd02d1 U131 ( .A1(n195), .A2(n211), .ZN(n182) );
  nr02d1 U132 ( .A1(n141), .A2(n140), .ZN(n139) );
  inv0d1 U133 ( .I(n144), .ZN(n140) );
  inv0d1 U134 ( .I(n151), .ZN(n150) );
  inv0d1 U135 ( .I(n185), .ZN(n192) );
  inv0d1 U136 ( .I(n184), .ZN(n194) );
  inv0d1 U137 ( .I(n187), .ZN(n175) );
  nd02d1 U138 ( .A1(n183), .A2(n184), .ZN(n177) );
  inv0d1 U139 ( .I(n189), .ZN(n174) );
  inv0d1 U140 ( .I(n143), .ZN(n171) );
  inv0d1 U141 ( .I(n1), .ZN(n155) );
  nd04d0 U142 ( .A1(n166), .A2(n156), .A3(n153), .A4(n161), .ZN(n141) );
  inv0d1 U144 ( .I(n157), .ZN(n166) );
  nd02d1 U145 ( .A1(n167), .A2(n164), .ZN(n147) );
  nd02d1 U146 ( .A1(n170), .A2(n165), .ZN(n153) );
  nd02d1 U147 ( .A1(n139), .A2(n162), .ZN(N74) );
  nd02d1 U148 ( .A1(n139), .A2(n163), .ZN(N72) );
  inv0d1 U149 ( .I(n149), .ZN(n148) );
  nd02d1 U151 ( .A1(n181), .A2(n184), .ZN(n188) );
  nd02d1 U152 ( .A1(n181), .A2(n182), .ZN(n179) );
  inv0d1 U153 ( .I(pm66en), .ZN(n198) );
  inv0d1 U154 ( .I(pperr_n_in), .ZN(n204) );
  inv0d1 U155 ( .I(pidsel), .ZN(n209) );
  inv0d1 U156 ( .I(pserr_n_in), .ZN(n210) );
  an04d1 U157 ( .A1(pc_be_in[2]), .A2(pc_be_in[0]), .A3(n137), .A4(n138), .Z(
        n135) );
  an04d1 U158 ( .A1(pc_be_in[2]), .A2(pc_be_in[3]), .A3(n136), .A4(n137), .Z(
        n134) );
  nd02d1 U159 ( .A1(n201), .A2(n202), .ZN(n184) );
  nr04d0 U162 ( .A1(n138), .A2(n137), .A3(pc_be_in[0]), .A4(pc_be_in[2]), .ZN(
        n130) );
  nr04d0 U163 ( .A1(n137), .A2(n136), .A3(pc_be_in[2]), .A4(pc_be_in[3]), .ZN(
        n131) );
  nd02d1 U164 ( .A1(pstop_n_in), .A2(ppar_in), .ZN(n187) );
  inv0d1 U166 ( .I(pc_be_in[1]), .ZN(n137) );
  inv0d1 U167 ( .I(pgnt_n), .ZN(n207) );
  inv0d1 U169 ( .I(pframe_n_in), .ZN(n206) );
  inv0d1 U170 ( .I(pdevsel_n_in), .ZN(n203) );
  inv0d1 U171 ( .I(ptrdy_n_in), .ZN(n205) );
  inv0d1 U175 ( .I(pc_be_in[3]), .ZN(n138) );
  inv0d1 U176 ( .I(pc_be_in[0]), .ZN(n136) );
  inv0d1 U177 ( .I(pirdy_n_in), .ZN(n197) );
  nd02d1 U178 ( .A1(write_data[12]), .A2(n139), .ZN(n146) );
  nd02d1 U179 ( .A1(write_data[0]), .A2(n139), .ZN(n160) );
  nd02d1 U180 ( .A1(write_data[6]), .A2(n139), .ZN(n152) );
  inv0d1 U181 ( .I(write_empty), .ZN(n154) );
  inv0d1 U182 ( .I(cmd_in_valid), .ZN(n165) );
  bufbd1 U215 ( .I(cmd_in[1]), .Z(n1) );
  bufbd1 U218 ( .I(cmd_in[1]), .Z(n214) );
  inv0d1 U242 ( .I(cmd_in[3]), .ZN(n169) );
  inv0d1 U244 ( .I(cmd_in[0]), .ZN(n163) );
  inv0d1 U293 ( .I(cmd_in[2]), .ZN(n162) );
  oaim211d1 U294 ( .C1(write_data[14]), .C2(n139), .A(n144), .B(n145), .ZN(N90) );
endmodule


module SD_W_MUX ( blender_data, pci_read_data, risc_result_data, sd_w_select, 
        sd_wfifo_data );
  input [31:0] blender_data;
  input [31:0] pci_read_data;
  input [31:0] risc_result_data;
  input [1:0] sd_w_select;
  output [31:0] sd_wfifo_data;
  wire   n3, n4, n5, n6, n1, n2, n7, n8, n9, n10, n11, n12, n13;

  an02d1 U1 ( .A1(sd_w_select[0]), .A2(n6), .Z(n5) );
  aor222d1 U3 ( .A1(risc_result_data[9]), .A2(n13), .B1(pci_read_data[9]), 
        .B2(n8), .C1(blender_data[9]), .C2(n1), .Z(sd_wfifo_data[9]) );
  aor222d1 U4 ( .A1(risc_result_data[8]), .A2(n13), .B1(pci_read_data[8]), 
        .B2(n8), .C1(blender_data[8]), .C2(n1), .Z(sd_wfifo_data[8]) );
  aor222d1 U5 ( .A1(risc_result_data[7]), .A2(n13), .B1(pci_read_data[7]), 
        .B2(n8), .C1(blender_data[7]), .C2(n1), .Z(sd_wfifo_data[7]) );
  aor222d1 U6 ( .A1(risc_result_data[6]), .A2(n13), .B1(pci_read_data[6]), 
        .B2(n8), .C1(blender_data[6]), .C2(n1), .Z(sd_wfifo_data[6]) );
  aor222d1 U7 ( .A1(risc_result_data[5]), .A2(n13), .B1(pci_read_data[5]), 
        .B2(n8), .C1(blender_data[5]), .C2(n1), .Z(sd_wfifo_data[5]) );
  aor222d1 U8 ( .A1(risc_result_data[4]), .A2(n13), .B1(pci_read_data[4]), 
        .B2(n8), .C1(blender_data[4]), .C2(n1), .Z(sd_wfifo_data[4]) );
  aor222d1 U9 ( .A1(risc_result_data[3]), .A2(n13), .B1(pci_read_data[3]), 
        .B2(n8), .C1(blender_data[3]), .C2(n1), .Z(sd_wfifo_data[3]) );
  aor222d1 U10 ( .A1(risc_result_data[31]), .A2(n13), .B1(pci_read_data[31]), 
        .B2(n8), .C1(blender_data[31]), .C2(n1), .Z(sd_wfifo_data[31]) );
  aor222d1 U11 ( .A1(risc_result_data[30]), .A2(n12), .B1(pci_read_data[30]), 
        .B2(n8), .C1(blender_data[30]), .C2(n1), .Z(sd_wfifo_data[30]) );
  aor222d1 U12 ( .A1(risc_result_data[2]), .A2(n12), .B1(pci_read_data[2]), 
        .B2(n8), .C1(blender_data[2]), .C2(n1), .Z(sd_wfifo_data[2]) );
  aor222d1 U13 ( .A1(risc_result_data[29]), .A2(n12), .B1(pci_read_data[29]), 
        .B2(n8), .C1(blender_data[29]), .C2(n1), .Z(sd_wfifo_data[29]) );
  aor222d1 U14 ( .A1(risc_result_data[28]), .A2(n12), .B1(pci_read_data[28]), 
        .B2(n8), .C1(blender_data[28]), .C2(n1), .Z(sd_wfifo_data[28]) );
  aor222d1 U15 ( .A1(risc_result_data[27]), .A2(n12), .B1(pci_read_data[27]), 
        .B2(n9), .C1(blender_data[27]), .C2(n2), .Z(sd_wfifo_data[27]) );
  aor222d1 U16 ( .A1(risc_result_data[26]), .A2(n12), .B1(pci_read_data[26]), 
        .B2(n9), .C1(blender_data[26]), .C2(n2), .Z(sd_wfifo_data[26]) );
  aor222d1 U17 ( .A1(risc_result_data[25]), .A2(n12), .B1(pci_read_data[25]), 
        .B2(n9), .C1(blender_data[25]), .C2(n2), .Z(sd_wfifo_data[25]) );
  aor222d1 U18 ( .A1(risc_result_data[24]), .A2(n12), .B1(pci_read_data[24]), 
        .B2(n9), .C1(blender_data[24]), .C2(n2), .Z(sd_wfifo_data[24]) );
  aor222d1 U19 ( .A1(risc_result_data[23]), .A2(n12), .B1(pci_read_data[23]), 
        .B2(n9), .C1(blender_data[23]), .C2(n2), .Z(sd_wfifo_data[23]) );
  aor222d1 U20 ( .A1(risc_result_data[22]), .A2(n12), .B1(pci_read_data[22]), 
        .B2(n9), .C1(blender_data[22]), .C2(n2), .Z(sd_wfifo_data[22]) );
  aor222d1 U21 ( .A1(risc_result_data[21]), .A2(n12), .B1(pci_read_data[21]), 
        .B2(n9), .C1(blender_data[21]), .C2(n2), .Z(sd_wfifo_data[21]) );
  aor222d1 U22 ( .A1(risc_result_data[20]), .A2(n12), .B1(pci_read_data[20]), 
        .B2(n9), .C1(blender_data[20]), .C2(n2), .Z(sd_wfifo_data[20]) );
  aor222d1 U23 ( .A1(risc_result_data[1]), .A2(n11), .B1(pci_read_data[1]), 
        .B2(n9), .C1(blender_data[1]), .C2(n2), .Z(sd_wfifo_data[1]) );
  aor222d1 U24 ( .A1(risc_result_data[19]), .A2(n11), .B1(pci_read_data[19]), 
        .B2(n9), .C1(blender_data[19]), .C2(n2), .Z(sd_wfifo_data[19]) );
  aor222d1 U25 ( .A1(risc_result_data[18]), .A2(n11), .B1(pci_read_data[18]), 
        .B2(n9), .C1(blender_data[18]), .C2(n2), .Z(sd_wfifo_data[18]) );
  aor222d1 U26 ( .A1(risc_result_data[17]), .A2(n11), .B1(pci_read_data[17]), 
        .B2(n9), .C1(blender_data[17]), .C2(n2), .Z(sd_wfifo_data[17]) );
  aor222d1 U27 ( .A1(risc_result_data[16]), .A2(n11), .B1(pci_read_data[16]), 
        .B2(n10), .C1(blender_data[16]), .C2(n7), .Z(sd_wfifo_data[16]) );
  aor222d1 U28 ( .A1(risc_result_data[15]), .A2(n11), .B1(pci_read_data[15]), 
        .B2(n10), .C1(blender_data[15]), .C2(n7), .Z(sd_wfifo_data[15]) );
  aor222d1 U29 ( .A1(risc_result_data[14]), .A2(n11), .B1(pci_read_data[14]), 
        .B2(n10), .C1(blender_data[14]), .C2(n7), .Z(sd_wfifo_data[14]) );
  aor222d1 U30 ( .A1(risc_result_data[13]), .A2(n11), .B1(pci_read_data[13]), 
        .B2(n10), .C1(blender_data[13]), .C2(n7), .Z(sd_wfifo_data[13]) );
  aor222d1 U31 ( .A1(risc_result_data[12]), .A2(n11), .B1(pci_read_data[12]), 
        .B2(n10), .C1(blender_data[12]), .C2(n7), .Z(sd_wfifo_data[12]) );
  aor222d1 U32 ( .A1(risc_result_data[11]), .A2(n11), .B1(pci_read_data[11]), 
        .B2(n10), .C1(blender_data[11]), .C2(n7), .Z(sd_wfifo_data[11]) );
  aor222d1 U33 ( .A1(risc_result_data[10]), .A2(n11), .B1(pci_read_data[10]), 
        .B2(n10), .C1(blender_data[10]), .C2(n7), .Z(sd_wfifo_data[10]) );
  aor222d1 U34 ( .A1(risc_result_data[0]), .A2(n11), .B1(pci_read_data[0]), 
        .B2(n10), .C1(blender_data[0]), .C2(n7), .Z(sd_wfifo_data[0]) );
  xn02d1 U35 ( .A1(sd_w_select[0]), .A2(sd_w_select[1]), .ZN(n4) );
  nr02d0 U36 ( .A1(n6), .A2(sd_w_select[0]), .ZN(n3) );
  bufbd1 U2 ( .I(n3), .Z(n11) );
  bufbd1 U37 ( .I(n3), .Z(n12) );
  bufbd1 U38 ( .I(n5), .Z(n2) );
  bufbd1 U39 ( .I(n5), .Z(n1) );
  bufbd1 U40 ( .I(n4), .Z(n9) );
  bufbd1 U41 ( .I(n4), .Z(n8) );
  bufbd1 U42 ( .I(n3), .Z(n13) );
  bufbd1 U43 ( .I(n5), .Z(n7) );
  bufbd1 U44 ( .I(n4), .Z(n10) );
  inv0d1 U45 ( .I(sd_w_select[1]), .ZN(n6) );
endmodule


module PCI_W_MUX ( blender_data, sdram_read_data, risc_result_data, 
        pci_w_select, pci_wfifo_data );
  input [31:0] blender_data;
  input [31:0] sdram_read_data;
  input [31:0] risc_result_data;
  input [1:0] pci_w_select;
  output [31:0] pci_wfifo_data;
  wire   n3, n4, n5, n6, n1, n2, n7, n8, n9, n10, n11, n12, n13;

  an02d1 U1 ( .A1(pci_w_select[0]), .A2(n6), .Z(n5) );
  aor222d1 U3 ( .A1(sdram_read_data[9]), .A2(n13), .B1(risc_result_data[9]), 
        .B2(n8), .C1(blender_data[9]), .C2(n1), .Z(pci_wfifo_data[9]) );
  aor222d1 U4 ( .A1(sdram_read_data[8]), .A2(n13), .B1(risc_result_data[8]), 
        .B2(n8), .C1(blender_data[8]), .C2(n1), .Z(pci_wfifo_data[8]) );
  aor222d1 U5 ( .A1(sdram_read_data[7]), .A2(n13), .B1(risc_result_data[7]), 
        .B2(n8), .C1(blender_data[7]), .C2(n1), .Z(pci_wfifo_data[7]) );
  aor222d1 U6 ( .A1(sdram_read_data[6]), .A2(n13), .B1(risc_result_data[6]), 
        .B2(n8), .C1(blender_data[6]), .C2(n1), .Z(pci_wfifo_data[6]) );
  aor222d1 U7 ( .A1(sdram_read_data[5]), .A2(n13), .B1(risc_result_data[5]), 
        .B2(n8), .C1(blender_data[5]), .C2(n1), .Z(pci_wfifo_data[5]) );
  aor222d1 U8 ( .A1(sdram_read_data[4]), .A2(n13), .B1(risc_result_data[4]), 
        .B2(n8), .C1(blender_data[4]), .C2(n1), .Z(pci_wfifo_data[4]) );
  aor222d1 U9 ( .A1(sdram_read_data[3]), .A2(n13), .B1(risc_result_data[3]), 
        .B2(n8), .C1(blender_data[3]), .C2(n1), .Z(pci_wfifo_data[3]) );
  aor222d1 U10 ( .A1(sdram_read_data[31]), .A2(n13), .B1(risc_result_data[31]), 
        .B2(n8), .C1(blender_data[31]), .C2(n1), .Z(pci_wfifo_data[31]) );
  aor222d1 U11 ( .A1(sdram_read_data[30]), .A2(n12), .B1(risc_result_data[30]), 
        .B2(n8), .C1(blender_data[30]), .C2(n1), .Z(pci_wfifo_data[30]) );
  aor222d1 U12 ( .A1(sdram_read_data[2]), .A2(n12), .B1(risc_result_data[2]), 
        .B2(n8), .C1(blender_data[2]), .C2(n1), .Z(pci_wfifo_data[2]) );
  aor222d1 U13 ( .A1(sdram_read_data[29]), .A2(n12), .B1(risc_result_data[29]), 
        .B2(n8), .C1(blender_data[29]), .C2(n1), .Z(pci_wfifo_data[29]) );
  aor222d1 U14 ( .A1(sdram_read_data[28]), .A2(n12), .B1(risc_result_data[28]), 
        .B2(n8), .C1(blender_data[28]), .C2(n1), .Z(pci_wfifo_data[28]) );
  aor222d1 U15 ( .A1(sdram_read_data[27]), .A2(n12), .B1(risc_result_data[27]), 
        .B2(n9), .C1(blender_data[27]), .C2(n2), .Z(pci_wfifo_data[27]) );
  aor222d1 U16 ( .A1(sdram_read_data[26]), .A2(n12), .B1(risc_result_data[26]), 
        .B2(n9), .C1(blender_data[26]), .C2(n2), .Z(pci_wfifo_data[26]) );
  aor222d1 U17 ( .A1(sdram_read_data[25]), .A2(n12), .B1(risc_result_data[25]), 
        .B2(n9), .C1(blender_data[25]), .C2(n2), .Z(pci_wfifo_data[25]) );
  aor222d1 U18 ( .A1(sdram_read_data[24]), .A2(n12), .B1(risc_result_data[24]), 
        .B2(n9), .C1(blender_data[24]), .C2(n2), .Z(pci_wfifo_data[24]) );
  aor222d1 U19 ( .A1(sdram_read_data[23]), .A2(n12), .B1(risc_result_data[23]), 
        .B2(n9), .C1(blender_data[23]), .C2(n2), .Z(pci_wfifo_data[23]) );
  aor222d1 U20 ( .A1(sdram_read_data[22]), .A2(n12), .B1(risc_result_data[22]), 
        .B2(n9), .C1(blender_data[22]), .C2(n2), .Z(pci_wfifo_data[22]) );
  aor222d1 U21 ( .A1(sdram_read_data[21]), .A2(n12), .B1(risc_result_data[21]), 
        .B2(n9), .C1(blender_data[21]), .C2(n2), .Z(pci_wfifo_data[21]) );
  aor222d1 U22 ( .A1(sdram_read_data[20]), .A2(n12), .B1(risc_result_data[20]), 
        .B2(n9), .C1(blender_data[20]), .C2(n2), .Z(pci_wfifo_data[20]) );
  aor222d1 U23 ( .A1(sdram_read_data[1]), .A2(n11), .B1(risc_result_data[1]), 
        .B2(n9), .C1(blender_data[1]), .C2(n2), .Z(pci_wfifo_data[1]) );
  aor222d1 U24 ( .A1(sdram_read_data[19]), .A2(n11), .B1(risc_result_data[19]), 
        .B2(n9), .C1(blender_data[19]), .C2(n2), .Z(pci_wfifo_data[19]) );
  aor222d1 U25 ( .A1(sdram_read_data[18]), .A2(n11), .B1(risc_result_data[18]), 
        .B2(n9), .C1(blender_data[18]), .C2(n2), .Z(pci_wfifo_data[18]) );
  aor222d1 U26 ( .A1(sdram_read_data[17]), .A2(n11), .B1(risc_result_data[17]), 
        .B2(n9), .C1(blender_data[17]), .C2(n2), .Z(pci_wfifo_data[17]) );
  aor222d1 U27 ( .A1(sdram_read_data[16]), .A2(n11), .B1(risc_result_data[16]), 
        .B2(n10), .C1(blender_data[16]), .C2(n7), .Z(pci_wfifo_data[16]) );
  aor222d1 U28 ( .A1(sdram_read_data[15]), .A2(n11), .B1(risc_result_data[15]), 
        .B2(n10), .C1(blender_data[15]), .C2(n7), .Z(pci_wfifo_data[15]) );
  aor222d1 U29 ( .A1(sdram_read_data[14]), .A2(n11), .B1(risc_result_data[14]), 
        .B2(n10), .C1(blender_data[14]), .C2(n7), .Z(pci_wfifo_data[14]) );
  aor222d1 U30 ( .A1(sdram_read_data[13]), .A2(n11), .B1(risc_result_data[13]), 
        .B2(n10), .C1(blender_data[13]), .C2(n7), .Z(pci_wfifo_data[13]) );
  aor222d1 U31 ( .A1(sdram_read_data[12]), .A2(n11), .B1(risc_result_data[12]), 
        .B2(n10), .C1(blender_data[12]), .C2(n7), .Z(pci_wfifo_data[12]) );
  aor222d1 U32 ( .A1(sdram_read_data[11]), .A2(n11), .B1(risc_result_data[11]), 
        .B2(n10), .C1(blender_data[11]), .C2(n7), .Z(pci_wfifo_data[11]) );
  aor222d1 U33 ( .A1(sdram_read_data[10]), .A2(n11), .B1(risc_result_data[10]), 
        .B2(n10), .C1(blender_data[10]), .C2(n7), .Z(pci_wfifo_data[10]) );
  aor222d1 U34 ( .A1(sdram_read_data[0]), .A2(n11), .B1(risc_result_data[0]), 
        .B2(n10), .C1(blender_data[0]), .C2(n7), .Z(pci_wfifo_data[0]) );
  xn02d1 U35 ( .A1(pci_w_select[0]), .A2(pci_w_select[1]), .ZN(n4) );
  nr02d0 U36 ( .A1(n6), .A2(pci_w_select[0]), .ZN(n3) );
  bufbd1 U2 ( .I(n3), .Z(n11) );
  bufbd1 U37 ( .I(n3), .Z(n12) );
  bufbd1 U38 ( .I(n5), .Z(n2) );
  bufbd1 U39 ( .I(n5), .Z(n1) );
  bufbd1 U40 ( .I(n4), .Z(n9) );
  bufbd1 U41 ( .I(n4), .Z(n8) );
  bufbd1 U42 ( .I(n3), .Z(n13) );
  bufbd1 U43 ( .I(n5), .Z(n7) );
  bufbd1 U44 ( .I(n4), .Z(n10) );
  inv0d1 U45 ( .I(pci_w_select[1]), .ZN(n6) );
endmodule


module SDRAM_TOP ( sys_clk, sdram_clk, sys_rst_n, sdram_rst_n, test_mode, 
        risc_OUT_VALID, risc_STACK_FULL, risc_EndOfInstrn, risc_PSW, 
        risc_Rd_Instr, sd_A, sd_CK, sd_CKn, sd_LD, sd_RW, sd_BWS, sd_DQ_in, 
        sd_DQ_out, sd_DQ_en, sd_sys_data_out, sd_wfifo_data, 
        parser_sd_rfifo_pop, parser_sd_wfifo_push, sd_rfifo_parser_empty, 
        sd_wfifo_parser_full, test_si1, test_si2, test_si3, test_si4, test_si5, 
        test_se, test_so1, test_so3, test_so5 );
  input [10:0] risc_PSW;
  output [9:0] sd_A;
  output [1:0] sd_BWS;
  input [15:0] sd_DQ_in;
  output [15:0] sd_DQ_out;
  output [15:0] sd_DQ_en;
  output [31:0] sd_sys_data_out;
  input [31:0] sd_wfifo_data;
  input sys_clk, sdram_clk, sys_rst_n, sdram_rst_n, test_mode, risc_OUT_VALID,
         risc_STACK_FULL, risc_EndOfInstrn, risc_Rd_Instr, parser_sd_rfifo_pop,
         parser_sd_wfifo_push, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_se;
  output sd_CK, sd_CKn, sd_LD, sd_RW, sd_rfifo_parser_empty,
         sd_wfifo_parser_full, test_so1, test_so3, test_so5;
  wire   net_sd_wfifo_pop, net_sd_wfifo_empty, net_sd_rfifo_push,
         net_sd_rfifo_full, n3, n7, n9, n10, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40;
  wire   [31:0] net_sdram_if_rDQ;
  wire   [31:0] net_sdram_if_wDQ;

  SDRAM_IF I_SDRAM_IF ( .sdram_clk(sdram_clk), .sdram_rst_n(sdram_rst_n), 
        .risc_OUT_VALID(risc_OUT_VALID), .risc_STACK_FULL(risc_STACK_FULL), 
        .risc_EndOfInstrn(risc_EndOfInstrn), .risc_PSW(risc_PSW), 
        .risc_Rd_Instr(risc_Rd_Instr), .sd_A(sd_A), .sd_CK(sd_CK), .sd_CKn(
        sd_CKn), .sd_LD(sd_LD), .sd_RW(sd_RW), .sd_BWS(sd_BWS), .sd_DQ_in(
        sd_DQ_in), .sd_DQ_out(sd_DQ_out), .sd_DQ_en(sd_DQ_en), .sd_wfifo_pop(
        net_sd_wfifo_pop), .sd_wfifo_empty(net_sd_wfifo_empty), 
        .sd_rfifo_push(net_sd_rfifo_push), .sd_rfifo_full(net_sd_rfifo_full), 
        .sd_rfifo_DQ_out(net_sdram_if_rDQ), .sd_wfifo_DQ_in(net_sdram_if_wDQ), 
        .test_se(test_se), .test_si1(test_si2), .test_si2(test_si1), 
        .test_si3(n9), .test_so2(test_so1), .test_so1(n10) );
  SDRAM_FIFO_0 I_SDRAM_READ_FIFO ( .fifo_clk_push(sdram_clk), .fifo_clk_pop(
        sys_clk), .fifo_rst_n(sdram_rst_n), .test_mode(test_mode), 
        .fifo_push_req_n(net_sd_rfifo_push), .fifo_pop_req_n(
        parser_sd_rfifo_pop), .fifo_data_in(net_sdram_if_rDQ), 
        .push_empty_fifo(SYNOPSYS_UNCONNECTED_21), .push_ae_fifo(
        SYNOPSYS_UNCONNECTED_22), .push_hf_fifo(SYNOPSYS_UNCONNECTED_23), 
        .push_af_fifo(SYNOPSYS_UNCONNECTED_24), .push_full_fifo(
        net_sd_rfifo_full), .push_error_fifo(SYNOPSYS_UNCONNECTED_25), 
        .pop_empty_fifo(sd_rfifo_parser_empty), .pop_ae_fifo(
        SYNOPSYS_UNCONNECTED_26), .pop_hf_fifo(SYNOPSYS_UNCONNECTED_27), 
        .pop_af_fifo(SYNOPSYS_UNCONNECTED_28), .pop_full_fifo(
        SYNOPSYS_UNCONNECTED_29), .pop_error_fifo(SYNOPSYS_UNCONNECTED_30), 
        .data_out_fifo(sd_sys_data_out), .test_se(test_se), .test_si1(test_si5), .test_si2(n10), .test_si3(test_si4), .test_si4(test_si3), .test_so1(n3), 
        .test_so2(n9), .test_so4(n7) );
  SDRAM_FIFO_1 I_SDRAM_WRITE_FIFO ( .fifo_clk_push(sys_clk), .fifo_clk_pop(
        sdram_clk), .fifo_rst_n(sys_rst_n), .test_mode(test_mode), 
        .fifo_push_req_n(parser_sd_wfifo_push), .fifo_pop_req_n(
        net_sd_wfifo_pop), .fifo_data_in(sd_wfifo_data), .push_empty_fifo(
        SYNOPSYS_UNCONNECTED_31), .push_ae_fifo(SYNOPSYS_UNCONNECTED_32), 
        .push_hf_fifo(SYNOPSYS_UNCONNECTED_33), .push_af_fifo(
        SYNOPSYS_UNCONNECTED_34), .push_full_fifo(sd_wfifo_parser_full), 
        .push_error_fifo(SYNOPSYS_UNCONNECTED_35), .pop_empty_fifo(
        net_sd_wfifo_empty), .pop_ae_fifo(SYNOPSYS_UNCONNECTED_36), 
        .pop_hf_fifo(SYNOPSYS_UNCONNECTED_37), .pop_af_fifo(
        SYNOPSYS_UNCONNECTED_38), .pop_full_fifo(SYNOPSYS_UNCONNECTED_39), 
        .pop_error_fifo(SYNOPSYS_UNCONNECTED_40), .data_out_fifo(
        net_sdram_if_wDQ), .test_se(test_se), .test_si1(n7), .test_si2(n3), 
        .test_so1(test_so3), .test_so2(test_so5) );
endmodule


module BLENDER ( clk, reset_n, clk_enable, test_mode, operation, op1, op2, 
        result, test_se, test_si1, test_si2, test_so2, test_so1 );
  input [3:0] operation;
  input [31:0] op1;
  input [31:0] op2;
  output [31:0] result;
  input clk, reset_n, clk_enable, test_mode, test_se, test_si1, test_si2;
  output test_so2, test_so1;
  wire   latched_clk_en, gclk, trans1, trans2, trans3, rem_red, rem_blue,
         c_trans1, c_trans2, c_trans3, c_rem_red, c_rem_blue, c_rem_green,
         s1_op2_31_, s1_op2_30_, s1_op2_29_, s1_op2_28_, s1_op2_27_,
         s1_op2_26_, s1_op2_25_, s1_op2_24_, s1_op2_23_, s1_op2_22_,
         s1_op2_20_, s1_op2_19_, s1_op2_18_, s1_op2_17_, s1_op2_16_,
         s1_op2_15_, s1_op2_14_, s1_op2_13_, s1_op2_12_, s1_op2_11_,
         s1_op2_10_, s1_op2_9_, s1_op2_8_, s1_op2_7_, s1_op2_6_, s1_op2_5_,
         s1_op2_4_, s1_op2_3_, s1_op2_2_, s1_op2_1_, s1_op2_0_, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423,
         N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467,
         N468, N469, N470, N471, N472, N473, N474, N475, N476, N541, N542,
         N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564,
         N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575,
         N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597,
         N598, N599, N600, N601, N602, N603, N604, N607, N608, N609, N610,
         N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621,
         N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632,
         N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643,
         N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654,
         N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665,
         N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676,
         N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687,
         N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698,
         N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709,
         N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720,
         N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731,
         N732, N733, N734, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756,
         N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767,
         N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778,
         N779, N780, N781, N782, N783, N784, N785, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859,
         N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892,
         N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903,
         N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936,
         N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947,
         N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969,
         N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980,
         N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991,
         N992, N993, n440, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n469, n478, n479, n480,
         n481, n482, n484, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n468, n470, n471, n472, n473, n474, n475,
         n476, n477, n483, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16;
  wire   [31:0] s1_op1;
  wire   [31:0] s2_op1;
  wire   [31:0] s2_op2;
  wire   [31:0] s3_op1;
  wire   [31:0] s3_op2;
  wire   [31:0] s4_op1;
  wire   [31:0] s4_op2;
  wire   [15:0] s5_result;
  wire   [127:0] mega_shift;

  slnlq1 latched_clk_en_reg ( .D(clk_enable), .EN(clk), .SC(1'b0), .SD(n442), 
        .Q(latched_clk_en), .SO(n442) );
  sdcrn1 rem_green_reg ( .D(c_rem_green), .SD(rem_blue), .SC(test_se), .CP(
        gclk), .CDN(reset_n), .QN(n440) );
  or02d1 U451 ( .A1(c_rem_green), .A2(n461), .Z(c_trans2) );
  an02d1 U455 ( .A1(n459), .A2(operation[2]), .Z(c_rem_blue) );
  xr02d1 U467 ( .A1(s4_op2[19]), .A2(s4_op2[18]), .Z(n443) );
  xr02d1 U468 ( .A1(s4_op2[17]), .A2(s4_op2[16]), .Z(n444) );
  xr02d1 U469 ( .A1(s4_op2[15]), .A2(s4_op2[14]), .Z(n445) );
  xr02d1 U470 ( .A1(s4_op2[13]), .A2(s4_op2[12]), .Z(n446) );
  xr02d1 U471 ( .A1(s4_op2[11]), .A2(s4_op2[10]), .Z(n447) );
  xr02d1 U472 ( .A1(s4_op2[9]), .A2(s4_op2[8]), .Z(n448) );
  xr02d1 U473 ( .A1(s4_op2[7]), .A2(s4_op2[6]), .Z(n449) );
  xr02d1 U474 ( .A1(s4_op2[5]), .A2(s4_op2[4]), .Z(n450) );
  xr02d1 U475 ( .A1(s4_op2[3]), .A2(s4_op2[2]), .Z(n451) );
  xr02d1 U476 ( .A1(s4_op2[31]), .A2(s4_op2[30]), .Z(n452) );
  xr02d1 U477 ( .A1(s4_op2[29]), .A2(s4_op2[28]), .Z(n453) );
  xr02d1 U478 ( .A1(s4_op2[27]), .A2(s4_op2[26]), .Z(n454) );
  xr02d1 U479 ( .A1(s4_op2[25]), .A2(s4_op2[24]), .Z(n455) );
  xr02d1 U480 ( .A1(s4_op2[23]), .A2(s4_op2[22]), .Z(n456) );
  xr02d1 U481 ( .A1(s4_op2[21]), .A2(s4_op2[20]), .Z(n457) );
  xr02d1 U482 ( .A1(s4_op2[1]), .A2(s4_op2[0]), .Z(n458) );
  ora21d1 U483 ( .B1(latched_clk_en), .B2(test_mode), .A(clk), .Z(gclk) );
  aor21d1 U484 ( .B1(n459), .B2(n460), .A(n461), .Z(c_trans3) );
  nd04d0 U485 ( .A1(operation[2]), .A2(operation[0]), .A3(n463), .A4(n464), 
        .ZN(n462) );
  nr04d0 U486 ( .A1(n460), .A2(n463), .A3(n464), .A4(operation[0]), .ZN(n461)
         );
  nr03d0 U487 ( .A1(n465), .A2(n466), .A3(n460), .ZN(c_rem_red) );
  xr02d1 U488 ( .A1(operation[3]), .A2(operation[1]), .Z(n465) );
  nr04d0 U489 ( .A1(n463), .A2(n464), .A3(operation[0]), .A4(operation[2]), 
        .ZN(c_rem_green) );
  nr03d0 U490 ( .A1(n466), .A2(operation[1]), .A3(n464), .ZN(n459) );
  aor22d1 U491 ( .A1(op1[13]), .A2(n514), .B1(op2[21]), .B2(n507), .Z(N99) );
  aor22d1 U492 ( .A1(op1[12]), .A2(n514), .B1(op2[20]), .B2(n507), .Z(N98) );
  aor22d1 U493 ( .A1(op1[11]), .A2(n514), .B1(op2[19]), .B2(n507), .Z(N97) );
  aor22d1 U494 ( .A1(op1[10]), .A2(n514), .B1(op2[18]), .B2(n507), .Z(N96) );
  aor22d1 U495 ( .A1(op1[9]), .A2(n514), .B1(op2[17]), .B2(n507), .Z(N95) );
  aor22d1 U496 ( .A1(op1[8]), .A2(n514), .B1(op2[16]), .B2(n507), .Z(N94) );
  aor222d1 U497 ( .A1(op1[15]), .A2(n507), .B1(op1[7]), .B2(n496), .C1(n517), 
        .C2(op2[7]), .Z(N93) );
  aor222d1 U498 ( .A1(op1[14]), .A2(n507), .B1(op1[6]), .B2(n495), .C1(op2[6]), 
        .C2(n515), .Z(N92) );
  aor222d1 U499 ( .A1(op1[13]), .A2(n507), .B1(op1[5]), .B2(n469), .C1(op2[5]), 
        .C2(n515), .Z(N91) );
  aor222d1 U500 ( .A1(op1[12]), .A2(n506), .B1(op1[4]), .B2(n496), .C1(op2[4]), 
        .C2(n515), .Z(N90) );
  aor222d1 U509 ( .A1(op1[11]), .A2(n506), .B1(op1[3]), .B2(n495), .C1(op2[3]), 
        .C2(n515), .Z(N89) );
  aor222d1 U520 ( .A1(op1[10]), .A2(n506), .B1(op1[2]), .B2(n469), .C1(op2[2]), 
        .C2(n515), .Z(N88) );
  aor222d1 U531 ( .A1(op1[9]), .A2(n506), .B1(op1[1]), .B2(n496), .C1(op2[1]), 
        .C2(n515), .Z(N87) );
  aor222d1 U542 ( .A1(op1[8]), .A2(n506), .B1(op1[0]), .B2(n495), .C1(op2[0]), 
        .C2(n515), .Z(N86) );
  aor22d1 U636 ( .A1(s1_op1[7]), .A2(n498), .B1(s1_op2_31_), .B2(n479), .Z(
        N344) );
  aor22d1 U637 ( .A1(s1_op1[6]), .A2(n497), .B1(s1_op2_30_), .B2(n500), .Z(
        N343) );
  aor22d1 U638 ( .A1(s1_op1[5]), .A2(n478), .B1(s1_op2_29_), .B2(n499), .Z(
        N342) );
  aor22d1 U639 ( .A1(s1_op1[4]), .A2(n498), .B1(s1_op2_28_), .B2(n479), .Z(
        N341) );
  aor22d1 U640 ( .A1(s1_op1[3]), .A2(n497), .B1(s1_op2_27_), .B2(n500), .Z(
        N340) );
  aor22d1 U641 ( .A1(s1_op1[2]), .A2(n478), .B1(s1_op2_26_), .B2(n499), .Z(
        N339) );
  aor22d1 U642 ( .A1(s1_op1[1]), .A2(n498), .B1(s1_op2_25_), .B2(n479), .Z(
        N338) );
  aor22d1 U643 ( .A1(s1_op1[0]), .A2(n497), .B1(s1_op2_24_), .B2(n500), .Z(
        N337) );
  aor22d1 U644 ( .A1(s1_op1[23]), .A2(n501), .B1(s1_op2_23_), .B2(n499), .Z(
        N336) );
  aor22d1 U645 ( .A1(s1_op1[22]), .A2(n501), .B1(s1_op2_22_), .B2(n479), .Z(
        N335) );
  aor22d1 U646 ( .A1(s1_op1[21]), .A2(n501), .B1(test_so1), .B2(n500), .Z(N334) );
  aor22d1 U647 ( .A1(s1_op1[20]), .A2(n501), .B1(s1_op2_20_), .B2(n499), .Z(
        N333) );
  aor22d1 U648 ( .A1(s1_op1[19]), .A2(n501), .B1(s1_op2_19_), .B2(n479), .Z(
        N332) );
  aor22d1 U649 ( .A1(s1_op1[18]), .A2(n501), .B1(s1_op2_18_), .B2(n500), .Z(
        N331) );
  aor22d1 U650 ( .A1(s1_op1[17]), .A2(n501), .B1(s1_op2_17_), .B2(n499), .Z(
        N330) );
  aor22d1 U651 ( .A1(s1_op1[16]), .A2(n501), .B1(s1_op2_16_), .B2(n479), .Z(
        N329) );
  aor22d1 U652 ( .A1(s1_op2_15_), .A2(n481), .B1(n482), .B2(s1_op1[23]), .Z(
        N328) );
  aor22d1 U653 ( .A1(s1_op2_14_), .A2(n481), .B1(n482), .B2(s1_op1[22]), .Z(
        N327) );
  aor22d1 U654 ( .A1(s1_op2_13_), .A2(n481), .B1(n482), .B2(s1_op1[21]), .Z(
        N326) );
  aor22d1 U655 ( .A1(s1_op2_12_), .A2(n481), .B1(n482), .B2(s1_op1[20]), .Z(
        N325) );
  aor22d1 U656 ( .A1(s1_op2_11_), .A2(n481), .B1(n482), .B2(s1_op1[19]), .Z(
        N324) );
  aor22d1 U657 ( .A1(s1_op2_10_), .A2(n481), .B1(n482), .B2(s1_op1[18]), .Z(
        N323) );
  aor22d1 U658 ( .A1(s1_op2_9_), .A2(n481), .B1(n482), .B2(s1_op1[17]), .Z(
        N322) );
  aor22d1 U659 ( .A1(s1_op2_8_), .A2(n481), .B1(n482), .B2(s1_op1[16]), .Z(
        N321) );
  aor222d1 U660 ( .A1(s1_op2_15_), .A2(n478), .B1(s1_op2_7_), .B2(n500), .C1(
        s1_op1[7]), .C2(n492), .Z(N320) );
  aor222d1 U661 ( .A1(s1_op2_14_), .A2(n498), .B1(s1_op2_6_), .B2(n499), .C1(
        s1_op1[6]), .C2(n493), .Z(N319) );
  aor222d1 U662 ( .A1(s1_op2_13_), .A2(n497), .B1(s1_op2_5_), .B2(n479), .C1(
        s1_op1[5]), .C2(n492), .Z(N318) );
  aor222d1 U663 ( .A1(s1_op2_12_), .A2(n478), .B1(s1_op2_4_), .B2(n500), .C1(
        s1_op1[4]), .C2(n493), .Z(N317) );
  aor222d1 U664 ( .A1(s1_op2_11_), .A2(n498), .B1(s1_op2_3_), .B2(n499), .C1(
        s1_op1[3]), .C2(n494), .Z(N316) );
  aor222d1 U665 ( .A1(s1_op2_10_), .A2(n497), .B1(s1_op2_2_), .B2(n479), .C1(
        s1_op1[2]), .C2(n493), .Z(N315) );
  aor222d1 U666 ( .A1(s1_op2_9_), .A2(n478), .B1(s1_op2_1_), .B2(n500), .C1(
        s1_op1[1]), .C2(n494), .Z(N314) );
  aor222d1 U667 ( .A1(s1_op2_8_), .A2(n498), .B1(s1_op2_0_), .B2(n499), .C1(
        s1_op1[0]), .C2(n492), .Z(N313) );
  aor22d1 U668 ( .A1(s1_op2_7_), .A2(n497), .B1(s1_op1[31]), .B2(n479), .Z(
        N312) );
  aor22d1 U669 ( .A1(s1_op2_6_), .A2(n478), .B1(s1_op1[30]), .B2(n500), .Z(
        N311) );
  aor22d1 U670 ( .A1(s1_op2_5_), .A2(n498), .B1(s1_op1[29]), .B2(n499), .Z(
        N310) );
  aor22d1 U671 ( .A1(s1_op2_4_), .A2(n497), .B1(s1_op1[28]), .B2(n479), .Z(
        N309) );
  aor22d1 U672 ( .A1(s1_op2_3_), .A2(n478), .B1(s1_op1[27]), .B2(n500), .Z(
        N308) );
  aor22d1 U673 ( .A1(s1_op2_2_), .A2(n498), .B1(s1_op1[26]), .B2(n499), .Z(
        N307) );
  aor22d1 U674 ( .A1(s1_op2_1_), .A2(n497), .B1(s1_op1[25]), .B2(n479), .Z(
        N306) );
  aor22d1 U675 ( .A1(s1_op2_0_), .A2(n478), .B1(s1_op1[24]), .B2(n500), .Z(
        N305) );
  aor22d1 U676 ( .A1(s1_op2_23_), .A2(n501), .B1(s1_op1[23]), .B2(n499), .Z(
        N304) );
  aor22d1 U677 ( .A1(s1_op2_22_), .A2(n501), .B1(s1_op1[22]), .B2(n479), .Z(
        N303) );
  aor22d1 U678 ( .A1(test_so1), .A2(n501), .B1(s1_op1[21]), .B2(n500), .Z(N302) );
  aor22d1 U679 ( .A1(s1_op2_20_), .A2(n501), .B1(s1_op1[20]), .B2(n499), .Z(
        N301) );
  aor22d1 U680 ( .A1(s1_op2_19_), .A2(n501), .B1(s1_op1[19]), .B2(n479), .Z(
        N300) );
  aor22d1 U681 ( .A1(s1_op2_18_), .A2(n501), .B1(s1_op1[18]), .B2(n500), .Z(
        N299) );
  aor22d1 U682 ( .A1(s1_op2_17_), .A2(n501), .B1(s1_op1[17]), .B2(n499), .Z(
        N298) );
  aor22d1 U683 ( .A1(s1_op2_16_), .A2(n501), .B1(s1_op1[16]), .B2(n479), .Z(
        N297) );
  aor21d1 U684 ( .B1(rem_blue), .B2(n440), .A(n493), .Z(n480) );
  aor22d1 U685 ( .A1(s1_op1[15]), .A2(n481), .B1(n482), .B2(s1_op2_23_), .Z(
        N296) );
  aor22d1 U686 ( .A1(s1_op1[14]), .A2(n481), .B1(n482), .B2(s1_op2_22_), .Z(
        N295) );
  aor22d1 U687 ( .A1(s1_op1[13]), .A2(n481), .B1(n482), .B2(test_so1), .Z(N294) );
  aor22d1 U688 ( .A1(s1_op1[12]), .A2(n481), .B1(n482), .B2(s1_op2_20_), .Z(
        N293) );
  aor22d1 U689 ( .A1(s1_op1[11]), .A2(n481), .B1(n482), .B2(s1_op2_19_), .Z(
        N292) );
  aor22d1 U690 ( .A1(s1_op1[10]), .A2(n481), .B1(n482), .B2(s1_op2_18_), .Z(
        N291) );
  aor22d1 U691 ( .A1(s1_op1[9]), .A2(n481), .B1(n482), .B2(s1_op2_17_), .Z(
        N290) );
  aor22d1 U692 ( .A1(s1_op1[8]), .A2(n481), .B1(n482), .B2(s1_op2_16_), .Z(
        N289) );
  aor222d1 U694 ( .A1(s1_op1[15]), .A2(n498), .B1(s1_op1[7]), .B2(n500), .C1(
        s1_op2_7_), .C2(n494), .Z(N288) );
  aor222d1 U695 ( .A1(s1_op1[14]), .A2(n497), .B1(s1_op1[6]), .B2(n499), .C1(
        s1_op2_6_), .C2(n492), .Z(N287) );
  aor222d1 U696 ( .A1(s1_op1[13]), .A2(n498), .B1(s1_op1[5]), .B2(n479), .C1(
        s1_op2_5_), .C2(n493), .Z(N286) );
  aor222d1 U697 ( .A1(s1_op1[12]), .A2(n498), .B1(s1_op1[4]), .B2(n500), .C1(
        s1_op2_4_), .C2(n492), .Z(N285) );
  aor222d1 U698 ( .A1(s1_op1[11]), .A2(n497), .B1(s1_op1[3]), .B2(n499), .C1(
        s1_op2_3_), .C2(n493), .Z(N284) );
  aor222d1 U699 ( .A1(s1_op1[10]), .A2(n497), .B1(s1_op1[2]), .B2(n479), .C1(
        s1_op2_2_), .C2(n494), .Z(N283) );
  aor222d1 U700 ( .A1(s1_op1[9]), .A2(n498), .B1(s1_op1[1]), .B2(n500), .C1(
        s1_op2_1_), .C2(n493), .Z(N282) );
  aor222d1 U701 ( .A1(s1_op1[8]), .A2(n497), .B1(s1_op1[0]), .B2(n499), .C1(
        s1_op2_0_), .C2(n494), .Z(N281) );
  nr02d0 U704 ( .A1(n946), .A2(rem_blue), .ZN(n484) );
  aor22d1 U705 ( .A1(op2[31]), .A2(n514), .B1(op1[7]), .B2(n506), .Z(N149) );
  aor22d1 U706 ( .A1(op2[30]), .A2(n514), .B1(op1[6]), .B2(n506), .Z(N148) );
  aor22d1 U707 ( .A1(op2[29]), .A2(n513), .B1(op1[5]), .B2(n506), .Z(N147) );
  aor22d1 U708 ( .A1(op2[28]), .A2(n513), .B1(op1[4]), .B2(n506), .Z(N146) );
  aor22d1 U709 ( .A1(op2[27]), .A2(n513), .B1(op1[3]), .B2(n506), .Z(N145) );
  aor22d1 U710 ( .A1(op2[26]), .A2(n513), .B1(op1[2]), .B2(n506), .Z(N144) );
  aor22d1 U711 ( .A1(op2[25]), .A2(n512), .B1(op1[1]), .B2(n505), .Z(N143) );
  aor22d1 U712 ( .A1(op2[24]), .A2(n512), .B1(op1[0]), .B2(n505), .Z(N142) );
  aor222d1 U713 ( .A1(op2[31]), .A2(n505), .B1(op2[23]), .B2(n469), .C1(
        op1[23]), .C2(n515), .Z(N141) );
  aor222d1 U714 ( .A1(op2[30]), .A2(n505), .B1(op2[22]), .B2(n496), .C1(
        op1[22]), .C2(n515), .Z(N140) );
  aor222d1 U715 ( .A1(op2[29]), .A2(n505), .B1(n495), .B2(op2[21]), .C1(
        op1[21]), .C2(n515), .Z(N139) );
  aor222d1 U716 ( .A1(op2[28]), .A2(n505), .B1(n469), .B2(op2[20]), .C1(
        op1[20]), .C2(n515), .Z(N138) );
  aor222d1 U717 ( .A1(op2[27]), .A2(n505), .B1(n496), .B2(op2[19]), .C1(
        op1[19]), .C2(n515), .Z(N137) );
  aor222d1 U718 ( .A1(op2[26]), .A2(n505), .B1(n495), .B2(op2[18]), .C1(
        op1[18]), .C2(n515), .Z(N136) );
  aor222d1 U719 ( .A1(op2[25]), .A2(n505), .B1(n469), .B2(op2[17]), .C1(
        op1[17]), .C2(n515), .Z(N135) );
  aor222d1 U720 ( .A1(op2[24]), .A2(n505), .B1(n496), .B2(op2[16]), .C1(
        op1[16]), .C2(n516), .Z(N134) );
  aor22d1 U721 ( .A1(op2[15]), .A2(n512), .B1(op1[23]), .B2(n505), .Z(N133) );
  aor22d1 U722 ( .A1(op2[14]), .A2(n512), .B1(op1[22]), .B2(n504), .Z(N132) );
  aor22d1 U723 ( .A1(op2[13]), .A2(n511), .B1(op1[21]), .B2(n504), .Z(N131) );
  aor22d1 U724 ( .A1(op2[12]), .A2(n511), .B1(op1[20]), .B2(n504), .Z(N130) );
  aor22d1 U725 ( .A1(op2[11]), .A2(n511), .B1(op1[19]), .B2(n504), .Z(N129) );
  aor22d1 U726 ( .A1(op2[10]), .A2(n511), .B1(op1[18]), .B2(n504), .Z(N128) );
  aor22d1 U727 ( .A1(op2[9]), .A2(n510), .B1(op1[17]), .B2(n504), .Z(N127) );
  aor22d1 U728 ( .A1(op2[8]), .A2(n510), .B1(op1[16]), .B2(n504), .Z(N126) );
  aor222d1 U729 ( .A1(op2[15]), .A2(n504), .B1(op2[7]), .B2(n495), .C1(n516), 
        .C2(op1[7]), .Z(N125) );
  aor222d1 U730 ( .A1(op2[14]), .A2(n504), .B1(op2[6]), .B2(n469), .C1(op1[6]), 
        .C2(n516), .Z(N124) );
  aor222d1 U731 ( .A1(op2[13]), .A2(n504), .B1(op2[5]), .B2(n496), .C1(op1[5]), 
        .C2(n516), .Z(N123) );
  aor222d1 U732 ( .A1(op2[12]), .A2(n504), .B1(op2[4]), .B2(n495), .C1(op1[4]), 
        .C2(n516), .Z(N122) );
  aor222d1 U733 ( .A1(op2[11]), .A2(n503), .B1(op2[3]), .B2(n469), .C1(op1[3]), 
        .C2(n516), .Z(N121) );
  aor222d1 U734 ( .A1(op2[10]), .A2(n503), .B1(op2[2]), .B2(n496), .C1(op1[2]), 
        .C2(n516), .Z(N120) );
  aor222d1 U735 ( .A1(op2[9]), .A2(n503), .B1(op2[1]), .B2(n495), .C1(op1[1]), 
        .C2(n516), .Z(N119) );
  aor222d1 U736 ( .A1(op2[8]), .A2(n503), .B1(op2[0]), .B2(n469), .C1(op1[0]), 
        .C2(n516), .Z(N118) );
  aor22d1 U737 ( .A1(op1[31]), .A2(n510), .B1(op2[7]), .B2(n503), .Z(N117) );
  aor22d1 U738 ( .A1(op1[30]), .A2(n510), .B1(op2[6]), .B2(n503), .Z(N116) );
  aor22d1 U739 ( .A1(op1[29]), .A2(n509), .B1(op2[5]), .B2(n503), .Z(N115) );
  aor22d1 U740 ( .A1(op1[28]), .A2(n509), .B1(op2[4]), .B2(n503), .Z(N114) );
  aor22d1 U741 ( .A1(op1[27]), .A2(n509), .B1(op2[3]), .B2(n503), .Z(N113) );
  aor22d1 U742 ( .A1(op1[26]), .A2(n509), .B1(op2[2]), .B2(n503), .Z(N112) );
  aor22d1 U743 ( .A1(op1[25]), .A2(n508), .B1(op2[1]), .B2(n503), .Z(N111) );
  aor22d1 U744 ( .A1(op1[24]), .A2(n508), .B1(op2[0]), .B2(n502), .Z(N110) );
  aor222d1 U745 ( .A1(op1[31]), .A2(n502), .B1(op1[23]), .B2(n496), .C1(
        op2[23]), .C2(n516), .Z(N109) );
  aor222d1 U746 ( .A1(op1[30]), .A2(n502), .B1(op1[22]), .B2(n495), .C1(
        op2[22]), .C2(n516), .Z(N108) );
  aor222d1 U747 ( .A1(op1[29]), .A2(n502), .B1(op1[21]), .B2(n469), .C1(n516), 
        .C2(op2[21]), .Z(N107) );
  aor222d1 U748 ( .A1(op1[28]), .A2(n502), .B1(op1[20]), .B2(n496), .C1(n516), 
        .C2(op2[20]), .Z(N106) );
  aor222d1 U749 ( .A1(op1[27]), .A2(n502), .B1(op1[19]), .B2(n495), .C1(n516), 
        .C2(op2[19]), .Z(N105) );
  aor222d1 U750 ( .A1(op1[26]), .A2(n502), .B1(op1[18]), .B2(n469), .C1(n516), 
        .C2(op2[18]), .Z(N104) );
  aor222d1 U751 ( .A1(op1[25]), .A2(n502), .B1(op1[17]), .B2(n496), .C1(n516), 
        .C2(op2[17]), .Z(N103) );
  aor222d1 U752 ( .A1(op1[24]), .A2(n502), .B1(op1[16]), .B2(n495), .C1(n517), 
        .C2(op2[16]), .Z(N102) );
  aor22d1 U754 ( .A1(op1[15]), .A2(n508), .B1(op2[23]), .B2(n502), .Z(N101) );
  aor22d1 U755 ( .A1(op1[14]), .A2(n508), .B1(op2[22]), .B2(n502), .Z(N100) );
  BLENDER_DW_mult_uns_4 mult_174 ( .a(s3_op2[31:20]), .b(s3_op2[19:8]), 
        .product({N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, 
        N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, 
        N763, N762}) );
  BLENDER_DW_mult_uns_3 mult_173 ( .a(s3_op1[31:20]), .b(s3_op1[19:8]), 
        .product({N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, 
        N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, 
        N739, N738}) );
  BLENDER_DW_mult_uns_5 mult_50_L43980_C203 ( .a(mega_shift[95:80]), .b(
        mega_shift[79:64]), .product({N929, N928, N927, N926, N925, N924, N923, 
        N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, 
        N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, 
        N898}) );
  BLENDER_DW_mult_uns_6 mult_50_L43980_C203_I2 ( .a(mega_shift[63:48]), .b(
        mega_shift[47:32]), .product({N961, N960, N959, N958, N957, N956, N955, 
        N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, 
        N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, 
        N930}) );
  BLENDER_DW_mult_uns_9 mult_50_L43980_C203_I3 ( .a(mega_shift[31:16]), .b(
        mega_shift[15:0]), .product({N993, N992, N991, N990, N989, N988, N987, 
        N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, 
        N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, 
        N962}) );
  BLENDER_DW01_add_6 add_157 ( .A(s2_op1), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b1, 1'b0}), .CI(1'b0), .SUM({N444, N443, N442, N441, N440, 
        N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, 
        N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, 
        N415, N414, N413}), .CO(SYNOPSYS_UNCONNECTED_9) );
  BLENDER_DW01_sub_6 sub_158 ( .A(s2_op2), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b1}), .CI(1'b0), .DIFF({N476, N475, N474, N473, N472, 
        N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, 
        N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, 
        N447, N446, N445}), .CO(SYNOPSYS_UNCONNECTED_10) );
  BLENDER_DW01_sub_7 sub_155 ( .A(s2_op2), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b1, 1'b1}), .CI(1'b0), .DIFF({N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, 
        N380, N379, N378}), .CO(SYNOPSYS_UNCONNECTED_11) );
  BLENDER_DW01_add_7 add_154 ( .A(s2_op1), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1, 1'b1}), .CI(1'b0), .SUM({N377, N376, N375, N374, N373, 
        N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, 
        N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, 
        N348, N347, N346}), .CO(SYNOPSYS_UNCONNECTED_12) );
  BLENDER_DW01_add_0 add_170 ( .A(s3_op1[31:16]), .B(s3_op1[15:0]), .CI(1'b0), 
        .SUM({N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, 
        N611, N610, N609, N608, N607}), .CO(SYNOPSYS_UNCONNECTED_13) );
  BLENDER_DW01_add_1 add_171 ( .A(s3_op2[31:16]), .B(s3_op1[15:0]), .CI(1'b0), 
        .SUM({N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671}), .CO(SYNOPSYS_UNCONNECTED_14) );
  BLENDER_DW01_sub_0 sub_170 ( .A(s3_op2[31:16]), .B(s3_op2[15:0]), .CI(1'b0), 
        .DIFF({N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, 
        N628, N627, N626, N625, N624, N623}), .CO(SYNOPSYS_UNCONNECTED_15) );
  BLENDER_DW01_sub_1 sub_171 ( .A(s3_op2[31:16]), .B(s3_op1[15:0]), .CI(1'b0), 
        .DIFF({N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        N692, N691, N690, N689, N688, N687}), .CO(SYNOPSYS_UNCONNECTED_16) );
  BLENDER_DW_mult_uns_0 mult_170 ( .a({N622, N621, N620, N619, N618, N617, 
        N616, N615, N614, N613, N612, N611, N610, N609, N608, N607}), .b({N638, 
        N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, 
        N625, N624, N623}), .product({N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, 
        N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, 
        N639}) );
  BLENDER_DW_mult_uns_1 mult_171 ( .a({N686, N685, N684, N683, N682, N681, 
        N680, N679, N678, N677, N676, N675, N674, N673, N672, N671}), .b({N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, 
        N689, N688, N687}), .product({N734, N733, N732, N731, N730, N729, N728, 
        N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, 
        N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, 
        N703}) );
  sdnrq1 s4_op1_reg_31_ ( .D(N865), .SD(s4_op1[30]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[31]) );
  sdnrq1 s4_op1_reg_29_ ( .D(N863), .SD(s4_op1[28]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[29]) );
  sdnrq1 s4_op1_reg_27_ ( .D(N861), .SD(s4_op1[26]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[27]) );
  sdnrq1 s4_op1_reg_25_ ( .D(N859), .SD(s4_op1[24]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[25]) );
  sdnrq1 s4_op1_reg_23_ ( .D(N857), .SD(s4_op1[22]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[23]) );
  sdnrq1 s4_op1_reg_21_ ( .D(N855), .SD(s4_op1[20]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[21]) );
  sdnrq1 s4_op1_reg_19_ ( .D(N853), .SD(s4_op1[18]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[19]) );
  sdnrq1 s4_op1_reg_17_ ( .D(N851), .SD(s4_op1[16]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[17]) );
  sdnrq1 s4_op1_reg_15_ ( .D(N849), .SD(s4_op1[14]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[15]) );
  sdnrq1 s4_op1_reg_13_ ( .D(N847), .SD(s4_op1[12]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[13]) );
  sdnrq1 s4_op1_reg_11_ ( .D(N845), .SD(s4_op1[10]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[11]) );
  sdnrq1 s4_op1_reg_9_ ( .D(N843), .SD(s4_op1[8]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[9]) );
  sdnrq1 s4_op1_reg_7_ ( .D(N841), .SD(s4_op1[6]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[7]) );
  sdnrq1 s4_op1_reg_5_ ( .D(N839), .SD(s4_op1[4]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[5]) );
  sdnrq1 s4_op1_reg_3_ ( .D(N837), .SD(s4_op1[2]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[3]) );
  sdnrq1 s4_op1_reg_1_ ( .D(N835), .SD(s4_op1[0]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[1]) );
  sdnrq1 s1_op2_reg_31_ ( .D(N149), .SD(s1_op2_30_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_31_) );
  sdnrq1 s1_op2_reg_30_ ( .D(N148), .SD(s1_op2_29_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_30_) );
  sdnrq1 s1_op2_reg_29_ ( .D(N147), .SD(s1_op2_28_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_29_) );
  sdnrq1 s1_op2_reg_28_ ( .D(N146), .SD(s1_op2_27_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_28_) );
  sdnrq1 s1_op2_reg_27_ ( .D(N145), .SD(s1_op2_26_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_27_) );
  sdnrq1 s1_op2_reg_26_ ( .D(N144), .SD(s1_op2_25_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_26_) );
  sdnrq1 s1_op2_reg_25_ ( .D(N143), .SD(s1_op2_24_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_25_) );
  sdnrq1 s1_op2_reg_24_ ( .D(N142), .SD(s1_op2_23_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_24_) );
  sdnrq1 s1_op1_reg_31_ ( .D(N117), .SD(s1_op1[30]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[31]) );
  sdnrq1 s1_op1_reg_30_ ( .D(N116), .SD(s1_op1[29]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[30]) );
  sdnrq1 s1_op1_reg_29_ ( .D(N115), .SD(s1_op1[28]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[29]) );
  sdnrq1 s1_op1_reg_28_ ( .D(N114), .SD(s1_op1[27]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[28]) );
  sdnrq1 s1_op1_reg_27_ ( .D(N113), .SD(s1_op1[26]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[27]) );
  sdnrq1 s1_op1_reg_26_ ( .D(N112), .SD(s1_op1[25]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[26]) );
  sdnrq1 s1_op1_reg_25_ ( .D(N111), .SD(s1_op1[24]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[25]) );
  sdnrq1 s1_op1_reg_24_ ( .D(N110), .SD(s1_op1[23]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[24]) );
  sdnrq1 s1_op2_reg_15_ ( .D(N133), .SD(s1_op2_14_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_15_) );
  sdnrq1 s1_op2_reg_14_ ( .D(N132), .SD(s1_op2_13_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_14_) );
  sdnrq1 s1_op2_reg_13_ ( .D(N131), .SD(s1_op2_12_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_13_) );
  sdnrq1 s1_op2_reg_12_ ( .D(N130), .SD(s1_op2_11_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_12_) );
  sdnrq1 s1_op2_reg_11_ ( .D(N129), .SD(s1_op2_10_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_11_) );
  sdnrq1 s1_op2_reg_10_ ( .D(N128), .SD(s1_op2_9_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_10_) );
  sdnrq1 s1_op2_reg_9_ ( .D(N127), .SD(s1_op2_8_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_9_) );
  sdnrq1 s1_op2_reg_8_ ( .D(N126), .SD(s1_op2_7_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_8_) );
  sdnrq1 s1_op1_reg_15_ ( .D(N101), .SD(s1_op1[14]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[15]) );
  sdnrq1 s1_op1_reg_14_ ( .D(N100), .SD(s1_op1[13]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[14]) );
  sdnrq1 s1_op1_reg_13_ ( .D(N99), .SD(s1_op1[12]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[13]) );
  sdnrq1 s1_op1_reg_12_ ( .D(N98), .SD(s1_op1[11]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[12]) );
  sdnrq1 s1_op1_reg_11_ ( .D(N97), .SD(s1_op1[10]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[11]) );
  sdnrq1 s1_op1_reg_10_ ( .D(N96), .SD(s1_op1[9]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[10]) );
  sdnrq1 s1_op1_reg_9_ ( .D(N95), .SD(s1_op1[8]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[9]) );
  sdnrq1 s1_op1_reg_8_ ( .D(N94), .SD(s1_op1[7]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[8]) );
  sdnrq1 s1_op2_reg_23_ ( .D(N141), .SD(s1_op2_22_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_23_) );
  sdnrq1 s1_op2_reg_22_ ( .D(N140), .SD(test_si2), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_22_) );
  sdnrq1 s1_op2_reg_21_ ( .D(N139), .SD(s1_op2_20_), .SC(test_se), .CP(gclk), 
        .Q(test_so1) );
  sdnrq1 s1_op2_reg_20_ ( .D(N138), .SD(s1_op2_19_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_20_) );
  sdnrq1 s1_op2_reg_19_ ( .D(N137), .SD(s1_op2_18_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_19_) );
  sdnrq1 s1_op2_reg_18_ ( .D(N136), .SD(s1_op2_17_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_18_) );
  sdnrq1 s1_op2_reg_17_ ( .D(N135), .SD(s1_op2_16_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_17_) );
  sdnrq1 s1_op2_reg_16_ ( .D(N134), .SD(s1_op2_15_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_16_) );
  sdnrq1 s1_op1_reg_23_ ( .D(N109), .SD(s1_op1[22]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[23]) );
  sdnrq1 s1_op1_reg_22_ ( .D(N108), .SD(s1_op1[21]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[22]) );
  sdnrq1 s1_op1_reg_21_ ( .D(N107), .SD(s1_op1[20]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[21]) );
  sdnrq1 s1_op1_reg_20_ ( .D(N106), .SD(s1_op1[19]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[20]) );
  sdnrq1 s1_op1_reg_19_ ( .D(N105), .SD(s1_op1[18]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[19]) );
  sdnrq1 s1_op1_reg_18_ ( .D(N104), .SD(s1_op1[17]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[18]) );
  sdnrq1 s1_op1_reg_17_ ( .D(N103), .SD(s1_op1[16]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[17]) );
  sdnrq1 s1_op1_reg_16_ ( .D(N102), .SD(s1_op1[15]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[16]) );
  sdnrq1 s4_op2_reg_30_ ( .D(N896), .SD(s4_op2[29]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[30]) );
  sdnrq1 s4_op2_reg_28_ ( .D(N894), .SD(s4_op2[27]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[28]) );
  sdnrq1 s4_op2_reg_26_ ( .D(N892), .SD(s4_op2[25]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[26]) );
  sdnrq1 s4_op2_reg_24_ ( .D(N890), .SD(s4_op2[23]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[24]) );
  sdnrq1 s4_op2_reg_22_ ( .D(N888), .SD(s4_op2[21]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[22]) );
  sdnrq1 s4_op2_reg_20_ ( .D(N886), .SD(s4_op2[19]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[20]) );
  sdnrq1 s4_op2_reg_18_ ( .D(N884), .SD(s4_op2[17]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[18]) );
  sdnrq1 s4_op2_reg_16_ ( .D(N882), .SD(s4_op2[15]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[16]) );
  sdnrq1 s4_op2_reg_14_ ( .D(N880), .SD(s4_op2[13]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[14]) );
  sdnrq1 s4_op2_reg_12_ ( .D(N878), .SD(s4_op2[11]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[12]) );
  sdnrq1 s4_op2_reg_10_ ( .D(N876), .SD(s4_op2[9]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[10]) );
  sdnrq1 s4_op2_reg_8_ ( .D(N874), .SD(s4_op2[7]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[8]) );
  sdnrq1 s4_op2_reg_6_ ( .D(N872), .SD(s4_op2[5]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[6]) );
  sdnrq1 s4_op2_reg_4_ ( .D(N870), .SD(s4_op2[3]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[4]) );
  sdnrq1 s4_op2_reg_2_ ( .D(N868), .SD(s4_op2[1]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[2]) );
  sdnrq1 s4_op2_reg_0_ ( .D(N866), .SD(s4_op1[31]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[0]) );
  sdnrq1 s4_op2_reg_31_ ( .D(N897), .SD(s4_op2[30]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[31]) );
  sdnrq1 s4_op2_reg_29_ ( .D(N895), .SD(s4_op2[28]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[29]) );
  sdnrq1 s4_op2_reg_27_ ( .D(N893), .SD(s4_op2[26]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[27]) );
  sdnrq1 s4_op2_reg_25_ ( .D(N891), .SD(s4_op2[24]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[25]) );
  sdnrq1 s4_op2_reg_23_ ( .D(N889), .SD(s4_op2[22]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[23]) );
  sdnrq1 s4_op2_reg_21_ ( .D(N887), .SD(s4_op2[20]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[21]) );
  sdnrq1 s4_op2_reg_19_ ( .D(N885), .SD(s4_op2[18]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[19]) );
  sdnrq1 s4_op2_reg_17_ ( .D(N883), .SD(s4_op2[16]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[17]) );
  sdnrq1 s4_op2_reg_15_ ( .D(N881), .SD(s4_op2[14]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[15]) );
  sdnrq1 s4_op2_reg_13_ ( .D(N879), .SD(s4_op2[12]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[13]) );
  sdnrq1 s4_op2_reg_11_ ( .D(N877), .SD(s4_op2[10]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[11]) );
  sdnrq1 s4_op2_reg_9_ ( .D(N875), .SD(s4_op2[8]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[9]) );
  sdnrq1 s4_op2_reg_7_ ( .D(N873), .SD(s4_op2[6]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[7]) );
  sdnrq1 s4_op2_reg_5_ ( .D(N871), .SD(s4_op2[4]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[5]) );
  sdnrq1 s4_op2_reg_3_ ( .D(N869), .SD(s4_op2[2]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[3]) );
  sdnrq1 s4_op2_reg_1_ ( .D(N867), .SD(s4_op2[0]), .SC(test_se), .CP(gclk), 
        .Q(s4_op2[1]) );
  sdnrq1 s4_op1_reg_30_ ( .D(N864), .SD(s4_op1[29]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[30]) );
  sdnrq1 s4_op1_reg_28_ ( .D(N862), .SD(s4_op1[27]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[28]) );
  sdnrq1 s4_op1_reg_26_ ( .D(N860), .SD(s4_op1[25]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[26]) );
  sdnrq1 s4_op1_reg_24_ ( .D(N858), .SD(s4_op1[23]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[24]) );
  sdnrq1 s4_op1_reg_22_ ( .D(N856), .SD(s4_op1[21]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[22]) );
  sdnrq1 s4_op1_reg_20_ ( .D(N854), .SD(s4_op1[19]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[20]) );
  sdnrq1 s4_op1_reg_18_ ( .D(N852), .SD(s4_op1[17]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[18]) );
  sdnrq1 s4_op1_reg_16_ ( .D(N850), .SD(s4_op1[15]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[16]) );
  sdnrq1 s4_op1_reg_14_ ( .D(N848), .SD(s4_op1[13]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[14]) );
  sdnrq1 s4_op1_reg_12_ ( .D(N846), .SD(s4_op1[11]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[12]) );
  sdnrq1 s4_op1_reg_10_ ( .D(N844), .SD(s4_op1[9]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[10]) );
  sdnrq1 s4_op1_reg_8_ ( .D(N842), .SD(s4_op1[7]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[8]) );
  sdnrq1 s4_op1_reg_6_ ( .D(N840), .SD(s4_op1[5]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[6]) );
  sdnrq1 s4_op1_reg_4_ ( .D(N838), .SD(s4_op1[3]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[4]) );
  sdnrq1 s4_op1_reg_2_ ( .D(N836), .SD(s4_op1[1]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[2]) );
  sdnrq1 s4_op1_reg_0_ ( .D(N834), .SD(s3_op2[31]), .SC(test_se), .CP(gclk), 
        .Q(s4_op1[0]) );
  sdcrq1 rem_blue_reg ( .D(c_rem_blue), .SD(mega_shift[31]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(rem_blue) );
  sdcrq1 result_reg_31_ ( .D(mega_shift[127]), .SD(result[30]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[31]) );
  sdcrq1 result_reg_30_ ( .D(mega_shift[126]), .SD(result[29]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[30]) );
  sdcrq1 result_reg_29_ ( .D(mega_shift[125]), .SD(result[28]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[29]) );
  sdcrq1 result_reg_28_ ( .D(mega_shift[124]), .SD(result[27]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[28]) );
  sdcrq1 result_reg_27_ ( .D(mega_shift[123]), .SD(result[26]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[27]) );
  sdcrq1 result_reg_26_ ( .D(mega_shift[122]), .SD(result[25]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[26]) );
  sdcrq1 result_reg_25_ ( .D(mega_shift[121]), .SD(result[24]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[25]) );
  sdcrq1 result_reg_24_ ( .D(mega_shift[120]), .SD(result[23]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[24]) );
  sdcrq1 result_reg_23_ ( .D(mega_shift[119]), .SD(result[22]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[23]) );
  sdcrq1 result_reg_22_ ( .D(mega_shift[118]), .SD(result[21]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[22]) );
  sdcrq1 result_reg_21_ ( .D(mega_shift[117]), .SD(result[20]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[21]) );
  sdcrq1 result_reg_20_ ( .D(mega_shift[116]), .SD(result[19]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[20]) );
  sdcrq1 result_reg_19_ ( .D(mega_shift[115]), .SD(result[18]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[19]) );
  sdcrq1 result_reg_18_ ( .D(mega_shift[114]), .SD(result[17]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[18]) );
  sdcrq1 result_reg_17_ ( .D(mega_shift[113]), .SD(result[16]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[17]) );
  sdcrq1 result_reg_16_ ( .D(mega_shift[112]), .SD(result[15]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[16]) );
  sdcrq1 result_reg_15_ ( .D(mega_shift[111]), .SD(result[14]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[15]) );
  sdcrq1 result_reg_14_ ( .D(mega_shift[110]), .SD(result[13]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[14]) );
  sdcrq1 result_reg_13_ ( .D(mega_shift[109]), .SD(result[12]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[13]) );
  sdcrq1 result_reg_12_ ( .D(mega_shift[108]), .SD(result[11]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[12]) );
  sdcrq1 result_reg_11_ ( .D(mega_shift[107]), .SD(result[10]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[11]) );
  sdcrq1 result_reg_10_ ( .D(mega_shift[106]), .SD(result[9]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[10]) );
  sdcrq1 result_reg_9_ ( .D(mega_shift[105]), .SD(result[8]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[9]) );
  sdcrq1 result_reg_8_ ( .D(mega_shift[104]), .SD(result[7]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[8]) );
  sdcrq1 result_reg_7_ ( .D(mega_shift[103]), .SD(result[6]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[7]) );
  sdcrq1 result_reg_6_ ( .D(mega_shift[102]), .SD(result[5]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[6]) );
  sdcrq1 result_reg_5_ ( .D(mega_shift[101]), .SD(result[4]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[5]) );
  sdcrq1 result_reg_4_ ( .D(mega_shift[100]), .SD(result[3]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[4]) );
  sdcrq1 result_reg_3_ ( .D(mega_shift[99]), .SD(result[2]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[3]) );
  sdcrq1 result_reg_2_ ( .D(mega_shift[98]), .SD(result[1]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[2]) );
  sdcrq1 result_reg_1_ ( .D(mega_shift[97]), .SD(result[0]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(result[1]) );
  sdcrq1 result_reg_0_ ( .D(mega_shift[96]), .SD(n493), .SC(test_se), .CP(gclk), .CDN(reset_n), .Q(result[0]) );
  sdnrq1 s1_op2_reg_7_ ( .D(N125), .SD(s1_op2_6_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_7_) );
  sdnrq1 s1_op2_reg_6_ ( .D(N124), .SD(s1_op2_5_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_6_) );
  sdnrq1 s1_op2_reg_5_ ( .D(N123), .SD(s1_op2_4_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_5_) );
  sdnrq1 s1_op2_reg_4_ ( .D(N122), .SD(s1_op2_3_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_4_) );
  sdnrq1 s1_op2_reg_3_ ( .D(N121), .SD(s1_op2_2_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_3_) );
  sdnrq1 s1_op2_reg_2_ ( .D(N120), .SD(s1_op2_1_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_2_) );
  sdnrq1 s1_op2_reg_1_ ( .D(N119), .SD(s1_op2_0_), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_1_) );
  sdnrq1 s1_op2_reg_0_ ( .D(N118), .SD(s1_op1[31]), .SC(test_se), .CP(gclk), 
        .Q(s1_op2_0_) );
  sdnrq1 s1_op1_reg_7_ ( .D(N93), .SD(s1_op1[6]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[7]) );
  sdnrq1 s1_op1_reg_6_ ( .D(N92), .SD(s1_op1[5]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[6]) );
  sdnrq1 s1_op1_reg_5_ ( .D(N91), .SD(s1_op1[4]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[5]) );
  sdnrq1 s1_op1_reg_4_ ( .D(N90), .SD(s1_op1[3]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[4]) );
  sdnrq1 s1_op1_reg_3_ ( .D(N89), .SD(s1_op1[2]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[3]) );
  sdnrq1 s1_op1_reg_2_ ( .D(N88), .SD(s1_op1[1]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[2]) );
  sdnrq1 s1_op1_reg_1_ ( .D(N87), .SD(s1_op1[0]), .SC(test_se), .CP(gclk), .Q(
        s1_op1[1]) );
  sdnrq1 s1_op1_reg_0_ ( .D(N86), .SD(result[31]), .SC(test_se), .CP(gclk), 
        .Q(s1_op1[0]) );
  sdnrq1 s2_op1_reg_31_ ( .D(N312), .SD(s2_op1[30]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[31]) );
  sdnrq1 s2_op2_reg_31_ ( .D(N344), .SD(s2_op2[30]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[31]) );
  sdnrq1 s2_op1_reg_30_ ( .D(N311), .SD(s2_op1[29]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[30]) );
  sdnrq1 s2_op1_reg_29_ ( .D(N310), .SD(s2_op1[28]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[29]) );
  sdnrq1 s2_op1_reg_28_ ( .D(N309), .SD(s2_op1[27]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[28]) );
  sdnrq1 s2_op1_reg_27_ ( .D(N308), .SD(s2_op1[26]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[27]) );
  sdcrq1 rem_red_reg ( .D(c_rem_red), .SD(n440), .SC(test_se), .CP(gclk), 
        .CDN(reset_n), .Q(rem_red) );
  sdcrq1 trans1_reg ( .D(c_trans1), .SD(s4_op2[31]), .SC(test_se), .CP(gclk), 
        .CDN(reset_n), .Q(trans1) );
  sdnrq1 s2_op2_reg_30_ ( .D(N343), .SD(s2_op2[29]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[30]) );
  sdnrq1 s2_op2_reg_29_ ( .D(N342), .SD(s2_op2[28]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[29]) );
  sdnrq1 s2_op2_reg_28_ ( .D(N341), .SD(s2_op2[27]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[28]) );
  sdnrq1 s2_op2_reg_27_ ( .D(N340), .SD(s2_op2[26]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[27]) );
  sdnrq1 s2_op2_reg_26_ ( .D(N339), .SD(s2_op2[25]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[26]) );
  sdcrq1 trans2_reg ( .D(c_trans2), .SD(n516), .SC(test_se), .CP(gclk), .CDN(
        reset_n), .Q(trans2) );
  sdcrq1 trans3_reg ( .D(c_trans3), .SD(trans2), .SC(test_se), .CP(gclk), 
        .CDN(reset_n), .Q(trans3) );
  sdnrq1 s2_op1_reg_26_ ( .D(N307), .SD(s2_op1[25]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[26]) );
  sdnrq1 s2_op1_reg_25_ ( .D(N306), .SD(s2_op1[24]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[25]) );
  sdnrq1 s2_op1_reg_24_ ( .D(N305), .SD(s2_op1[23]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[24]) );
  sdnrq1 s2_op1_reg_23_ ( .D(N304), .SD(s2_op1[22]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[23]) );
  sdnrq1 s2_op1_reg_22_ ( .D(N303), .SD(s2_op1[21]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[22]) );
  sdnrq1 s2_op1_reg_21_ ( .D(N302), .SD(s2_op1[20]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[21]) );
  sdnrq1 s2_op2_reg_25_ ( .D(N338), .SD(s2_op2[24]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[25]) );
  sdnrq1 s2_op2_reg_24_ ( .D(N337), .SD(s2_op2[23]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[24]) );
  sdnrq1 s2_op2_reg_23_ ( .D(N336), .SD(s2_op2[22]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[23]) );
  sdnrq1 s2_op2_reg_22_ ( .D(N335), .SD(s2_op2[21]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[22]) );
  sdnrq1 s2_op2_reg_21_ ( .D(N334), .SD(s2_op2[20]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[21]) );
  sdnrq1 s2_op2_reg_20_ ( .D(N333), .SD(s2_op2[19]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[20]) );
  sdnrq1 s2_op2_reg_19_ ( .D(N332), .SD(s2_op2[18]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[19]) );
  sdnrq1 s2_op1_reg_20_ ( .D(N301), .SD(s2_op1[19]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[20]) );
  sdnrq1 s2_op1_reg_19_ ( .D(N300), .SD(s2_op1[18]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[19]) );
  sdnrq1 s2_op1_reg_18_ ( .D(N299), .SD(s2_op1[17]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[18]) );
  sdnrq1 s2_op1_reg_17_ ( .D(N298), .SD(s2_op1[16]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[17]) );
  sdnrq1 s2_op1_reg_16_ ( .D(N297), .SD(s2_op1[15]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[16]) );
  sdnrq1 s2_op2_reg_18_ ( .D(N331), .SD(s2_op2[17]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[18]) );
  sdnrq1 s2_op2_reg_17_ ( .D(N330), .SD(s2_op2[16]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[17]) );
  sdnrq1 s2_op2_reg_16_ ( .D(N329), .SD(s2_op2[15]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[16]) );
  sdnrq1 s2_op2_reg_15_ ( .D(N328), .SD(s2_op2[14]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[15]) );
  sdnrq1 s2_op2_reg_14_ ( .D(N327), .SD(s2_op2[13]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[14]) );
  sdnrq1 s2_op2_reg_13_ ( .D(N326), .SD(s2_op2[12]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[13]) );
  sdnrq1 s2_op2_reg_12_ ( .D(N325), .SD(s2_op2[11]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[12]) );
  sdnrq1 s2_op1_reg_15_ ( .D(N296), .SD(s2_op1[14]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[15]) );
  sdnrq1 s2_op1_reg_14_ ( .D(N295), .SD(s2_op1[13]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[14]) );
  sdnrq1 s2_op1_reg_13_ ( .D(N294), .SD(s2_op1[12]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[13]) );
  sdnrq1 s2_op1_reg_12_ ( .D(N293), .SD(s2_op1[11]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[12]) );
  sdnrq1 s2_op1_reg_11_ ( .D(N292), .SD(s2_op1[10]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[11]) );
  sdnrq1 s2_op2_reg_9_ ( .D(N322), .SD(s2_op2[8]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[9]) );
  sdnrq1 s2_op2_reg_8_ ( .D(N321), .SD(s2_op2[7]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[8]) );
  sdnrq1 s2_op2_reg_11_ ( .D(N324), .SD(s2_op2[10]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[11]) );
  sdnrq1 s2_op2_reg_10_ ( .D(N323), .SD(s2_op2[9]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[10]) );
  sdnrq1 s2_op2_reg_7_ ( .D(N320), .SD(s2_op2[6]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[7]) );
  sdnrq1 s2_op2_reg_5_ ( .D(N318), .SD(s2_op2[4]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[5]) );
  sdnrq1 s2_op2_reg_4_ ( .D(N317), .SD(s2_op2[3]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[4]) );
  sdnrq1 s2_op2_reg_6_ ( .D(N319), .SD(s2_op2[5]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[6]) );
  sdnrq1 s2_op1_reg_10_ ( .D(N291), .SD(s2_op1[9]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[10]) );
  sdnrq1 s2_op1_reg_9_ ( .D(N290), .SD(s2_op1[8]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[9]) );
  sdnrq1 s2_op1_reg_8_ ( .D(N289), .SD(s2_op1[7]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[8]) );
  sdnrq1 s2_op2_reg_1_ ( .D(N314), .SD(s2_op2[0]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[1]) );
  sdnrq1 s2_op1_reg_0_ ( .D(N281), .SD(s1_op2_31_), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[0]) );
  sdnrq1 s2_op1_reg_5_ ( .D(N286), .SD(n761), .SC(test_se), .CP(gclk), .Q(
        s2_op1[5]) );
  sdnrq1 s2_op2_reg_2_ ( .D(N315), .SD(s2_op2[1]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[2]) );
  sdnrq1 s2_op1_reg_3_ ( .D(N284), .SD(n751), .SC(test_se), .CP(gclk), .Q(
        s2_op1[3]) );
  sdnrq1 s2_op1_reg_4_ ( .D(N285), .SD(n756), .SC(test_se), .CP(gclk), .Q(
        s2_op1[4]) );
  sdnrq1 s3_op1_reg_31_ ( .D(N572), .SD(s3_op1[30]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[31]) );
  sdnrq1 s2_op2_reg_3_ ( .D(N316), .SD(s2_op2[2]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[3]) );
  sdnrq1 s2_op1_reg_7_ ( .D(N288), .SD(s2_op1[6]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[7]) );
  sdnrq1 s2_op1_reg_6_ ( .D(N287), .SD(s2_op1[5]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[6]) );
  sdnrq1 s2_op2_reg_0_ ( .D(N313), .SD(s2_op1[31]), .SC(test_se), .CP(gclk), 
        .Q(s2_op2[0]) );
  sdnrq1 s3_op2_reg_31_ ( .D(N604), .SD(s3_op2[30]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[31]) );
  sdnrq1 s2_op1_reg_2_ ( .D(N283), .SD(n746), .SC(test_se), .CP(gclk), .Q(
        s2_op1[2]) );
  sdnrq1 s3_op2_reg_15_ ( .D(N588), .SD(n659), .SC(test_se), .CP(gclk), .Q(
        s3_op2[15]) );
  sdnrq1 s3_op2_reg_14_ ( .D(N587), .SD(n654), .SC(test_se), .CP(gclk), .Q(
        s3_op2[14]) );
  sdnrq1 s3_op2_reg_13_ ( .D(N586), .SD(n649), .SC(test_se), .CP(gclk), .Q(
        s3_op2[13]) );
  sdnrq1 s2_op1_reg_1_ ( .D(N282), .SD(s2_op1[0]), .SC(test_se), .CP(gclk), 
        .Q(s2_op1[1]) );
  sdnrq1 s3_op1_reg_30_ ( .D(N571), .SD(s3_op1[29]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[30]) );
  sdnrq1 s3_op1_reg_29_ ( .D(N570), .SD(s3_op1[28]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[29]) );
  sdnrq1 s3_op1_reg_28_ ( .D(N569), .SD(s3_op1[27]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[28]) );
  sdnrq1 s3_op1_reg_27_ ( .D(N568), .SD(n609), .SC(test_se), .CP(gclk), .Q(
        s3_op1[27]) );
  sdnrq1 s3_op1_reg_26_ ( .D(N567), .SD(n604), .SC(test_se), .CP(gclk), .Q(
        s3_op1[26]) );
  sdnrq1 s3_op1_reg_15_ ( .D(N556), .SD(n549), .SC(test_se), .CP(gclk), .Q(
        s3_op1[15]) );
  sdnrq1 s3_op2_reg_30_ ( .D(N603), .SD(s3_op2[29]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[30]) );
  sdnrq1 s3_op2_reg_29_ ( .D(N602), .SD(s3_op2[28]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[29]) );
  sdnrq1 s3_op2_reg_28_ ( .D(N601), .SD(s3_op2[27]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[28]) );
  sdnrq1 s3_op2_reg_27_ ( .D(N600), .SD(n719), .SC(test_se), .CP(gclk), .Q(
        s3_op2[27]) );
  sdnrq1 s3_op2_reg_26_ ( .D(N599), .SD(n714), .SC(test_se), .CP(gclk), .Q(
        s3_op2[26]) );
  sdnrq1 s3_op2_reg_7_ ( .D(N580), .SD(s3_op2[6]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[7]) );
  sdnrq1 s3_op2_reg_6_ ( .D(N579), .SD(s3_op2[5]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[6]) );
  sdnrq1 s3_op2_reg_5_ ( .D(N578), .SD(s3_op2[4]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[5]) );
  sdnrq1 s3_op2_reg_4_ ( .D(N577), .SD(s3_op2[3]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[4]) );
  sdnrq1 s3_op2_reg_3_ ( .D(N576), .SD(s3_op2[2]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[3]) );
  sdnrq1 s3_op2_reg_2_ ( .D(N575), .SD(s3_op2[1]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[2]) );
  sdnrq1 s3_op2_reg_1_ ( .D(N574), .SD(s3_op2[0]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[1]) );
  sdnrq1 s3_op2_reg_0_ ( .D(N573), .SD(s3_op1[31]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[0]) );
  sdcrq1 mega_shift_reg_1__31_ ( .D(N961), .SD(mega_shift[94]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[95]) );
  sdcrq1 mega_shift_reg_1__30_ ( .D(N960), .SD(mega_shift[93]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[94]) );
  sdcrq1 mega_shift_reg_1__29_ ( .D(N959), .SD(mega_shift[92]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[93]) );
  sdcrq1 mega_shift_reg_1__28_ ( .D(N958), .SD(mega_shift[91]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[92]) );
  sdcrq1 mega_shift_reg_1__27_ ( .D(N957), .SD(mega_shift[90]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[91]) );
  sdcrq1 mega_shift_reg_1__26_ ( .D(N956), .SD(mega_shift[89]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[90]) );
  sdcrq1 mega_shift_reg_1__25_ ( .D(N955), .SD(mega_shift[88]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[89]) );
  sdcrq1 mega_shift_reg_1__24_ ( .D(N954), .SD(mega_shift[87]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[88]) );
  sdcrq1 mega_shift_reg_1__23_ ( .D(N953), .SD(mega_shift[86]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[87]) );
  sdcrq1 mega_shift_reg_1__22_ ( .D(N952), .SD(mega_shift[85]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[86]) );
  sdcrq1 mega_shift_reg_1__21_ ( .D(N951), .SD(mega_shift[84]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[85]) );
  sdcrq1 mega_shift_reg_1__20_ ( .D(N950), .SD(mega_shift[83]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[84]) );
  sdcrq1 mega_shift_reg_1__19_ ( .D(N949), .SD(mega_shift[82]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[83]) );
  sdcrq1 mega_shift_reg_1__18_ ( .D(N948), .SD(mega_shift[81]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[82]) );
  sdcrq1 mega_shift_reg_1__17_ ( .D(N947), .SD(mega_shift[80]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[81]) );
  sdcrq1 mega_shift_reg_1__16_ ( .D(N946), .SD(mega_shift[79]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[80]) );
  sdcrq1 mega_shift_reg_1__15_ ( .D(N945), .SD(mega_shift[78]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[79]) );
  sdcrq1 mega_shift_reg_1__14_ ( .D(N944), .SD(mega_shift[77]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[78]) );
  sdcrq1 mega_shift_reg_1__13_ ( .D(N943), .SD(mega_shift[76]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[77]) );
  sdcrq1 mega_shift_reg_1__12_ ( .D(N942), .SD(mega_shift[75]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[76]) );
  sdcrq1 mega_shift_reg_1__11_ ( .D(N941), .SD(mega_shift[74]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[75]) );
  sdcrq1 mega_shift_reg_1__10_ ( .D(N940), .SD(mega_shift[73]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[74]) );
  sdcrq1 mega_shift_reg_1__9_ ( .D(N939), .SD(mega_shift[72]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[73]) );
  sdcrq1 mega_shift_reg_1__8_ ( .D(N938), .SD(mega_shift[71]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[72]) );
  sdcrq1 mega_shift_reg_1__7_ ( .D(N937), .SD(mega_shift[70]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[71]) );
  sdcrq1 mega_shift_reg_1__6_ ( .D(N936), .SD(mega_shift[69]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[70]) );
  sdcrq1 mega_shift_reg_1__5_ ( .D(N935), .SD(mega_shift[68]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[69]) );
  sdcrq1 mega_shift_reg_1__4_ ( .D(N934), .SD(mega_shift[67]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[68]) );
  sdcrq1 mega_shift_reg_1__3_ ( .D(N933), .SD(mega_shift[66]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[67]) );
  sdcrq1 mega_shift_reg_1__2_ ( .D(N932), .SD(mega_shift[65]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[66]) );
  sdcrq1 mega_shift_reg_1__1_ ( .D(N931), .SD(mega_shift[64]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[65]) );
  sdcrq1 mega_shift_reg_1__0_ ( .D(N930), .SD(mega_shift[127]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[64]) );
  sdcrq1 mega_shift_reg_2__31_ ( .D(N993), .SD(mega_shift[62]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[63]) );
  sdcrq1 mega_shift_reg_2__30_ ( .D(N992), .SD(mega_shift[61]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[62]) );
  sdcrq1 mega_shift_reg_2__29_ ( .D(N991), .SD(mega_shift[60]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[61]) );
  sdcrq1 mega_shift_reg_2__28_ ( .D(N990), .SD(mega_shift[59]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[60]) );
  sdcrq1 mega_shift_reg_2__27_ ( .D(N989), .SD(mega_shift[58]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[59]) );
  sdcrq1 mega_shift_reg_2__26_ ( .D(N988), .SD(mega_shift[57]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[58]) );
  sdcrq1 mega_shift_reg_2__25_ ( .D(N987), .SD(mega_shift[56]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[57]) );
  sdcrq1 mega_shift_reg_2__24_ ( .D(N986), .SD(mega_shift[55]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[56]) );
  sdcrq1 mega_shift_reg_2__23_ ( .D(N985), .SD(mega_shift[54]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[55]) );
  sdcrq1 mega_shift_reg_2__22_ ( .D(N984), .SD(mega_shift[53]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[54]) );
  sdcrq1 mega_shift_reg_2__21_ ( .D(N983), .SD(mega_shift[52]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[53]) );
  sdcrq1 mega_shift_reg_2__20_ ( .D(N982), .SD(mega_shift[51]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[52]) );
  sdcrq1 mega_shift_reg_2__19_ ( .D(N981), .SD(mega_shift[50]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[51]) );
  sdcrq1 mega_shift_reg_2__18_ ( .D(N980), .SD(mega_shift[49]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[50]) );
  sdcrq1 mega_shift_reg_2__17_ ( .D(N979), .SD(mega_shift[48]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[49]) );
  sdcrq1 mega_shift_reg_2__16_ ( .D(N978), .SD(mega_shift[47]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[48]) );
  sdcrq1 mega_shift_reg_2__15_ ( .D(N977), .SD(mega_shift[46]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[47]) );
  sdcrq1 mega_shift_reg_2__14_ ( .D(N976), .SD(mega_shift[45]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[46]) );
  sdcrq1 mega_shift_reg_2__13_ ( .D(N975), .SD(mega_shift[44]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[45]) );
  sdcrq1 mega_shift_reg_2__12_ ( .D(N974), .SD(mega_shift[43]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[44]) );
  sdcrq1 mega_shift_reg_2__11_ ( .D(N973), .SD(mega_shift[42]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[43]) );
  sdcrq1 mega_shift_reg_2__10_ ( .D(N972), .SD(mega_shift[41]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[42]) );
  sdcrq1 mega_shift_reg_2__9_ ( .D(N971), .SD(mega_shift[40]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[41]) );
  sdcrq1 mega_shift_reg_2__8_ ( .D(N970), .SD(mega_shift[39]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[40]) );
  sdcrq1 mega_shift_reg_2__7_ ( .D(N969), .SD(mega_shift[38]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[39]) );
  sdcrq1 mega_shift_reg_2__6_ ( .D(N968), .SD(mega_shift[37]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[38]) );
  sdcrq1 mega_shift_reg_2__5_ ( .D(N967), .SD(mega_shift[36]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[37]) );
  sdcrq1 mega_shift_reg_2__4_ ( .D(N966), .SD(mega_shift[35]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[36]) );
  sdcrq1 mega_shift_reg_2__3_ ( .D(N965), .SD(mega_shift[34]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[35]) );
  sdcrq1 mega_shift_reg_2__2_ ( .D(N964), .SD(mega_shift[33]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[34]) );
  sdcrq1 mega_shift_reg_2__1_ ( .D(N963), .SD(mega_shift[32]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[33]) );
  sdcrq1 mega_shift_reg_2__0_ ( .D(N962), .SD(mega_shift[95]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[32]) );
  sdcrq1 mega_shift_reg_3__31_ ( .D(s5_result[15]), .SD(mega_shift[30]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[31]) );
  sdcrq1 mega_shift_reg_3__30_ ( .D(s5_result[14]), .SD(mega_shift[29]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[30]) );
  sdcrq1 mega_shift_reg_3__29_ ( .D(s5_result[13]), .SD(mega_shift[28]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[29]) );
  sdcrq1 mega_shift_reg_3__28_ ( .D(s5_result[12]), .SD(mega_shift[27]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[28]) );
  sdcrq1 mega_shift_reg_3__27_ ( .D(s5_result[11]), .SD(mega_shift[26]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[27]) );
  sdcrq1 mega_shift_reg_3__26_ ( .D(s5_result[10]), .SD(mega_shift[25]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[26]) );
  sdcrq1 mega_shift_reg_3__25_ ( .D(s5_result[9]), .SD(mega_shift[24]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[25]) );
  sdcrq1 mega_shift_reg_3__24_ ( .D(s5_result[8]), .SD(mega_shift[23]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[24]) );
  sdcrq1 mega_shift_reg_3__23_ ( .D(s5_result[7]), .SD(mega_shift[22]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[23]) );
  sdcrq1 mega_shift_reg_3__22_ ( .D(s5_result[6]), .SD(mega_shift[21]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[22]) );
  sdcrq1 mega_shift_reg_3__21_ ( .D(s5_result[5]), .SD(mega_shift[20]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[21]) );
  sdcrq1 mega_shift_reg_3__20_ ( .D(s5_result[4]), .SD(mega_shift[19]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[20]) );
  sdcrq1 mega_shift_reg_3__19_ ( .D(s5_result[3]), .SD(mega_shift[18]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[19]) );
  sdcrq1 mega_shift_reg_3__18_ ( .D(s5_result[2]), .SD(mega_shift[17]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[18]) );
  sdcrq1 mega_shift_reg_3__17_ ( .D(s5_result[1]), .SD(mega_shift[16]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[17]) );
  sdcrq1 mega_shift_reg_3__16_ ( .D(s5_result[0]), .SD(mega_shift[15]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[16]) );
  sdcrq1 mega_shift_reg_3__15_ ( .D(s5_result[15]), .SD(mega_shift[14]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[15]) );
  sdcrq1 mega_shift_reg_3__14_ ( .D(s5_result[14]), .SD(mega_shift[13]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[14]) );
  sdcrq1 mega_shift_reg_3__13_ ( .D(s5_result[13]), .SD(mega_shift[12]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[13]) );
  sdcrq1 mega_shift_reg_3__12_ ( .D(s5_result[12]), .SD(mega_shift[11]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[12]) );
  sdcrq1 mega_shift_reg_3__11_ ( .D(s5_result[11]), .SD(mega_shift[10]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[11]) );
  sdcrq1 mega_shift_reg_3__10_ ( .D(s5_result[10]), .SD(mega_shift[9]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[10]) );
  sdcrq1 mega_shift_reg_3__9_ ( .D(s5_result[9]), .SD(mega_shift[8]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[9]) );
  sdcrq1 mega_shift_reg_3__8_ ( .D(s5_result[8]), .SD(mega_shift[7]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[8]) );
  sdcrq1 mega_shift_reg_3__7_ ( .D(s5_result[7]), .SD(mega_shift[6]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[7]) );
  sdcrq1 mega_shift_reg_3__6_ ( .D(s5_result[6]), .SD(mega_shift[5]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[6]) );
  sdcrq1 mega_shift_reg_3__5_ ( .D(s5_result[5]), .SD(mega_shift[4]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[5]) );
  sdcrq1 mega_shift_reg_3__4_ ( .D(s5_result[4]), .SD(mega_shift[3]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[4]) );
  sdcrq1 mega_shift_reg_3__3_ ( .D(s5_result[3]), .SD(mega_shift[2]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[3]) );
  sdcrq1 mega_shift_reg_3__2_ ( .D(s5_result[2]), .SD(mega_shift[1]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[2]) );
  sdcrq1 mega_shift_reg_3__1_ ( .D(s5_result[1]), .SD(mega_shift[0]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[1]) );
  sdcrq1 mega_shift_reg_3__0_ ( .D(s5_result[0]), .SD(mega_shift[63]), .SC(
        test_se), .CP(gclk), .CDN(reset_n), .Q(mega_shift[0]) );
  sdnrq1 s3_op2_reg_10_ ( .D(N583), .SD(n634), .SC(test_se), .CP(gclk), .Q(
        s3_op2[10]) );
  sdnrq1 s3_op1_reg_7_ ( .D(N548), .SD(s3_op1[6]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[7]) );
  sdnrq1 s3_op1_reg_4_ ( .D(N545), .SD(s3_op1[3]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[4]) );
  sdnrq1 s3_op1_reg_3_ ( .D(N544), .SD(s3_op1[2]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[3]) );
  sdnrq1 s3_op1_reg_2_ ( .D(N543), .SD(s3_op1[1]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[2]) );
  sdnrq1 s3_op1_reg_0_ ( .D(N541), .SD(s2_op2[31]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[0]) );
  sdnrq1 s3_op1_reg_6_ ( .D(N547), .SD(s3_op1[5]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[6]) );
  sdnrq1 s3_op1_reg_5_ ( .D(N546), .SD(s3_op1[4]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[5]) );
  sdnrq1 s3_op1_reg_1_ ( .D(N542), .SD(s3_op1[0]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[1]) );
  sdnrq1 s3_op1_reg_10_ ( .D(N551), .SD(n524), .SC(test_se), .CP(gclk), .Q(
        s3_op1[10]) );
  sdnrq1 s3_op2_reg_12_ ( .D(N585), .SD(n644), .SC(test_se), .CP(gclk), .Q(
        s3_op2[12]) );
  sdnrq1 s3_op2_reg_11_ ( .D(N584), .SD(n639), .SC(test_se), .CP(gclk), .Q(
        s3_op2[11]) );
  sdnrq1 s3_op2_reg_9_ ( .D(N582), .SD(n629), .SC(test_se), .CP(gclk), .Q(
        s3_op2[9]) );
  sdnrq1 s3_op2_reg_8_ ( .D(N581), .SD(s3_op2[7]), .SC(test_se), .CP(gclk), 
        .Q(s3_op2[8]) );
  sdnrq1 s3_op1_reg_22_ ( .D(N563), .SD(n584), .SC(test_se), .CP(gclk), .Q(
        s3_op1[22]) );
  sdnrq1 s3_op1_reg_21_ ( .D(N562), .SD(n579), .SC(test_se), .CP(gclk), .Q(
        s3_op1[21]) );
  sdnrq1 s3_op1_reg_17_ ( .D(N558), .SD(n559), .SC(test_se), .CP(gclk), .Q(
        s3_op1[17]) );
  sdnrq1 s3_op1_reg_25_ ( .D(N566), .SD(n599), .SC(test_se), .CP(gclk), .Q(
        s3_op1[25]) );
  sdnrq1 s3_op1_reg_24_ ( .D(N565), .SD(n594), .SC(test_se), .CP(gclk), .Q(
        s3_op1[24]) );
  sdnrq1 s3_op1_reg_23_ ( .D(N564), .SD(n589), .SC(test_se), .CP(gclk), .Q(
        s3_op1[23]) );
  sdnrq1 s3_op1_reg_20_ ( .D(N561), .SD(n574), .SC(test_se), .CP(gclk), .Q(
        s3_op1[20]) );
  sdnrq1 s3_op1_reg_19_ ( .D(N560), .SD(n569), .SC(test_se), .CP(gclk), .Q(
        s3_op1[19]) );
  sdnrq1 s3_op1_reg_18_ ( .D(N559), .SD(n564), .SC(test_se), .CP(gclk), .Q(
        s3_op1[18]) );
  sdnrq1 s3_op1_reg_16_ ( .D(N557), .SD(n554), .SC(test_se), .CP(gclk), .Q(
        s3_op1[16]) );
  sdnrq1 s3_op1_reg_9_ ( .D(N550), .SD(n518), .SC(test_se), .CP(gclk), .Q(
        s3_op1[9]) );
  sdnrq1 s3_op1_reg_8_ ( .D(N549), .SD(s3_op1[7]), .SC(test_se), .CP(gclk), 
        .Q(s3_op1[8]) );
  sdnrq1 s3_op2_reg_21_ ( .D(N594), .SD(n689), .SC(test_se), .CP(gclk), .Q(
        s3_op2[21]) );
  sdnrq1 s3_op2_reg_23_ ( .D(N596), .SD(n699), .SC(test_se), .CP(gclk), .Q(
        s3_op2[23]) );
  sdnrq1 s3_op2_reg_22_ ( .D(N595), .SD(n694), .SC(test_se), .CP(gclk), .Q(
        s3_op2[22]) );
  sdnrq1 s3_op2_reg_19_ ( .D(N592), .SD(n679), .SC(test_se), .CP(gclk), .Q(
        s3_op2[19]) );
  sdnrq1 s3_op2_reg_17_ ( .D(N590), .SD(n669), .SC(test_se), .CP(gclk), .Q(
        s3_op2[17]) );
  sdnrq1 s3_op2_reg_25_ ( .D(N598), .SD(n709), .SC(test_se), .CP(gclk), .Q(
        s3_op2[25]) );
  sdnrq1 s3_op2_reg_24_ ( .D(N597), .SD(n704), .SC(test_se), .CP(gclk), .Q(
        s3_op2[24]) );
  sdnrq1 s3_op2_reg_20_ ( .D(N593), .SD(n684), .SC(test_se), .CP(gclk), .Q(
        s3_op2[20]) );
  sdnrq1 s3_op2_reg_18_ ( .D(N591), .SD(n674), .SC(test_se), .CP(gclk), .Q(
        s3_op2[18]) );
  sdnrq1 s3_op1_reg_14_ ( .D(N555), .SD(n544), .SC(test_se), .CP(gclk), .Q(
        s3_op1[14]) );
  sdnrq1 s3_op1_reg_13_ ( .D(N554), .SD(n539), .SC(test_se), .CP(gclk), .Q(
        s3_op1[13]) );
  sdnrq1 s3_op1_reg_12_ ( .D(N553), .SD(n534), .SC(test_se), .CP(gclk), .Q(
        s3_op1[12]) );
  sdnrq1 s3_op1_reg_11_ ( .D(N552), .SD(n529), .SC(test_se), .CP(gclk), .Q(
        s3_op1[11]) );
  sdnrq1 s3_op2_reg_16_ ( .D(N589), .SD(n664), .SC(test_se), .CP(gclk), .Q(
        s3_op2[16]) );
  sdcrq1 mega_shift_reg_0__31_ ( .D(N929), .SD(mega_shift[126]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[127]) );
  sdcrq1 mega_shift_reg_0__30_ ( .D(N928), .SD(mega_shift[125]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[126]) );
  sdcrq1 mega_shift_reg_0__29_ ( .D(N927), .SD(mega_shift[124]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[125]) );
  sdcrq1 mega_shift_reg_0__28_ ( .D(N926), .SD(mega_shift[123]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[124]) );
  sdcrq1 mega_shift_reg_0__27_ ( .D(N925), .SD(mega_shift[122]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[123]) );
  sdcrq1 mega_shift_reg_0__26_ ( .D(N924), .SD(mega_shift[121]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[122]) );
  sdcrq1 mega_shift_reg_0__25_ ( .D(N923), .SD(mega_shift[120]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[121]) );
  sdcrq1 mega_shift_reg_0__24_ ( .D(N922), .SD(mega_shift[119]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[120]) );
  sdcrq1 mega_shift_reg_0__23_ ( .D(N921), .SD(mega_shift[118]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[119]) );
  sdcrq1 mega_shift_reg_0__22_ ( .D(N920), .SD(mega_shift[117]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[118]) );
  sdcrq1 mega_shift_reg_0__21_ ( .D(N919), .SD(mega_shift[116]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[117]) );
  sdcrq1 mega_shift_reg_0__20_ ( .D(N918), .SD(mega_shift[115]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[116]) );
  sdcrq1 mega_shift_reg_0__19_ ( .D(N917), .SD(mega_shift[114]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[115]) );
  sdcrq1 mega_shift_reg_0__18_ ( .D(N916), .SD(mega_shift[113]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[114]) );
  sdcrq1 mega_shift_reg_0__17_ ( .D(N915), .SD(mega_shift[112]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[113]) );
  sdcrq1 mega_shift_reg_0__16_ ( .D(N914), .SD(mega_shift[111]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[112]) );
  sdcrq1 mega_shift_reg_0__15_ ( .D(N913), .SD(mega_shift[110]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[111]) );
  sdcrq1 mega_shift_reg_0__14_ ( .D(N912), .SD(mega_shift[109]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[110]) );
  sdcrq1 mega_shift_reg_0__13_ ( .D(N911), .SD(mega_shift[108]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[109]) );
  sdcrq1 mega_shift_reg_0__12_ ( .D(N910), .SD(mega_shift[107]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[108]) );
  sdcrq1 mega_shift_reg_0__11_ ( .D(N909), .SD(mega_shift[106]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[107]) );
  sdcrq1 mega_shift_reg_0__10_ ( .D(N908), .SD(mega_shift[105]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[106]) );
  sdcrq1 mega_shift_reg_0__9_ ( .D(N907), .SD(mega_shift[104]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[105]) );
  sdcrq1 mega_shift_reg_0__8_ ( .D(N906), .SD(mega_shift[103]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[104]) );
  sdcrq1 mega_shift_reg_0__7_ ( .D(N905), .SD(mega_shift[102]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[103]) );
  sdcrq1 mega_shift_reg_0__6_ ( .D(N904), .SD(mega_shift[101]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[102]) );
  sdcrq1 mega_shift_reg_0__5_ ( .D(N903), .SD(mega_shift[100]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[101]) );
  sdcrq1 mega_shift_reg_0__4_ ( .D(N902), .SD(mega_shift[99]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[100]) );
  sdcrq1 mega_shift_reg_0__3_ ( .D(N901), .SD(mega_shift[98]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[99]) );
  sdcrq1 mega_shift_reg_0__2_ ( .D(N900), .SD(mega_shift[97]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[98]) );
  sdcrq1 mega_shift_reg_0__1_ ( .D(N899), .SD(mega_shift[96]), .SC(test_se), 
        .CP(gclk), .CDN(reset_n), .Q(mega_shift[97]) );
  sdcrq1 mega_shift_reg_0__0_ ( .D(N898), .SD(test_si1), .SC(test_se), .CP(
        gclk), .CDN(reset_n), .Q(mega_shift[96]) );
  nd12d0 U12 ( .A1(n13), .A2(N756), .ZN(n610) );
  nd12d0 U13 ( .A1(n13), .A2(N780), .ZN(n720) );
  nd12d0 U14 ( .A1(n736), .A2(N779), .ZN(n715) );
  nd12d0 U15 ( .A1(n736), .A2(N752), .ZN(n590) );
  nd12d0 U16 ( .A1(n736), .A2(N755), .ZN(n605) );
  nd12d0 U17 ( .A1(n736), .A2(N776), .ZN(n700) );
  nd12d0 U18 ( .A1(n13), .A2(N777), .ZN(n705) );
  nd12d0 U19 ( .A1(n13), .A2(N753), .ZN(n595) );
  nd12d0 U433 ( .A1(n14), .A2(N754), .ZN(n600) );
  nd12d0 U435 ( .A1(n14), .A2(N778), .ZN(n710) );
  nd12d0 U436 ( .A1(n14), .A2(N748), .ZN(n570) );
  nd12d0 U437 ( .A1(n736), .A2(N749), .ZN(n575) );
  nd12d0 U438 ( .A1(n13), .A2(N750), .ZN(n580) );
  nd12d0 U439 ( .A1(n14), .A2(N751), .ZN(n585) );
  nd12d0 U440 ( .A1(n14), .A2(N772), .ZN(n680) );
  nd12d0 U441 ( .A1(n736), .A2(N773), .ZN(n685) );
  nd12d0 U442 ( .A1(n13), .A2(N774), .ZN(n690) );
  nd12d0 U443 ( .A1(n14), .A2(N775), .ZN(n695) );
  nd12d0 U444 ( .A1(n13), .A2(N744), .ZN(n550) );
  nd12d0 U445 ( .A1(n14), .A2(N745), .ZN(n555) );
  nd12d0 U446 ( .A1(n736), .A2(N746), .ZN(n560) );
  nd12d0 U447 ( .A1(n13), .A2(N747), .ZN(n565) );
  nd12d0 U448 ( .A1(n13), .A2(N768), .ZN(n660) );
  nd12d0 U449 ( .A1(n14), .A2(N769), .ZN(n665) );
  nd12d0 U450 ( .A1(n736), .A2(N770), .ZN(n670) );
  nd12d0 U452 ( .A1(n13), .A2(N771), .ZN(n675) );
  nd12d0 U453 ( .A1(n14), .A2(N742), .ZN(n540) );
  nd12d0 U454 ( .A1(n736), .A2(N743), .ZN(n545) );
  nd12d0 U456 ( .A1(n14), .A2(N766), .ZN(n650) );
  nd12d0 U457 ( .A1(n736), .A2(N767), .ZN(n655) );
  nd12d0 U458 ( .A1(n13), .A2(N741), .ZN(n535) );
  nd12d0 U459 ( .A1(n13), .A2(N765), .ZN(n645) );
  inv0d1 U460 ( .I(n483), .ZN(n488) );
  inv0d1 U461 ( .I(n483), .ZN(n487) );
  inv0d1 U462 ( .I(n483), .ZN(n489) );
  inv0d1 U463 ( .I(n483), .ZN(n475) );
  inv0d1 U464 ( .I(n483), .ZN(n476) );
  inv0d1 U465 ( .I(n483), .ZN(n477) );
  inv0d1 U466 ( .I(n483), .ZN(n485) );
  inv0d1 U501 ( .I(n483), .ZN(n486) );
  inv0d1 U502 ( .I(n483), .ZN(n490) );
  inv0d1 U503 ( .I(n1), .ZN(n8) );
  inv0d1 U504 ( .I(n1), .ZN(n9) );
  inv0d1 U505 ( .I(n1), .ZN(n10) );
  inv0d1 U506 ( .I(n478), .ZN(n481) );
  inv0d1 U507 ( .I(n1), .ZN(n12) );
  inv0d1 U508 ( .I(n1), .ZN(n11) );
  nd12d0 U510 ( .A1(n736), .A2(N740), .ZN(n530) );
  nd12d0 U511 ( .A1(n14), .A2(N739), .ZN(n525) );
  nd12d0 U512 ( .A1(n14), .A2(N763), .ZN(n635) );
  nd12d0 U513 ( .A1(n736), .A2(N764), .ZN(n640) );
  inv0d1 U514 ( .I(n4), .ZN(n470) );
  inv0d1 U515 ( .I(n3), .ZN(n471) );
  inv0d1 U516 ( .I(n4), .ZN(n17) );
  inv0d1 U517 ( .I(n4), .ZN(n468) );
  inv0d1 U518 ( .I(n2), .ZN(n5) );
  inv0d1 U519 ( .I(n3), .ZN(n472) );
  inv0d1 U521 ( .I(n3), .ZN(n473) );
  inv0d1 U522 ( .I(n2), .ZN(n7) );
  inv0d1 U523 ( .I(n2), .ZN(n6) );
  inv0d1 U524 ( .I(n513), .ZN(n502) );
  inv0d1 U525 ( .I(n512), .ZN(n503) );
  inv0d1 U526 ( .I(n511), .ZN(n504) );
  inv0d1 U527 ( .I(n510), .ZN(n505) );
  inv0d1 U528 ( .I(n509), .ZN(n506) );
  inv0d1 U529 ( .I(n508), .ZN(n507) );
  nd12d0 U530 ( .A1(n718), .A2(n717), .ZN(N891) );
  nd12d0 U532 ( .A1(n716), .A2(n715), .ZN(n718) );
  nd12d0 U533 ( .A1(n5), .A2(N728), .ZN(n717) );
  nd12d0 U534 ( .A1(n608), .A2(n607), .ZN(N859) );
  nd12d0 U535 ( .A1(n606), .A2(n605), .ZN(n608) );
  nd12d0 U536 ( .A1(n7), .A2(N664), .ZN(n607) );
  nd12d0 U537 ( .A1(n673), .A2(n672), .ZN(N882) );
  nd12d0 U538 ( .A1(n671), .A2(n670), .ZN(n673) );
  nd12d0 U539 ( .A1(n5), .A2(N719), .ZN(n672) );
  nd12d0 U540 ( .A1(n678), .A2(n677), .ZN(N883) );
  nd12d0 U541 ( .A1(n676), .A2(n675), .ZN(n678) );
  nd12d0 U543 ( .A1(n5), .A2(N720), .ZN(n677) );
  nd12d0 U544 ( .A1(n683), .A2(n682), .ZN(N884) );
  nd12d0 U545 ( .A1(n681), .A2(n680), .ZN(n683) );
  nd12d0 U546 ( .A1(n5), .A2(N721), .ZN(n682) );
  nd12d0 U547 ( .A1(n688), .A2(n687), .ZN(N885) );
  nd12d0 U548 ( .A1(n686), .A2(n685), .ZN(n688) );
  nd12d0 U549 ( .A1(n5), .A2(N722), .ZN(n687) );
  nd12d0 U550 ( .A1(n693), .A2(n692), .ZN(N886) );
  nd12d0 U551 ( .A1(n691), .A2(n690), .ZN(n693) );
  nd12d0 U552 ( .A1(n5), .A2(N723), .ZN(n692) );
  nd12d0 U553 ( .A1(n698), .A2(n697), .ZN(N887) );
  nd12d0 U554 ( .A1(n696), .A2(n695), .ZN(n698) );
  nd12d0 U555 ( .A1(n5), .A2(N724), .ZN(n697) );
  nd12d0 U556 ( .A1(n713), .A2(n712), .ZN(N890) );
  nd12d0 U557 ( .A1(n711), .A2(n710), .ZN(n713) );
  nd12d0 U558 ( .A1(n5), .A2(N727), .ZN(n712) );
  nd12d0 U559 ( .A1(n723), .A2(n722), .ZN(N892) );
  nd12d0 U560 ( .A1(n721), .A2(n720), .ZN(n723) );
  nd12d0 U561 ( .A1(n5), .A2(N729), .ZN(n722) );
  nd12d0 U562 ( .A1(n563), .A2(n562), .ZN(N850) );
  nd12d0 U563 ( .A1(n561), .A2(n560), .ZN(n563) );
  nd12d0 U564 ( .A1(n6), .A2(N655), .ZN(n562) );
  nd12d0 U565 ( .A1(n568), .A2(n567), .ZN(N851) );
  nd12d0 U566 ( .A1(n566), .A2(n565), .ZN(n568) );
  nd12d0 U567 ( .A1(n7), .A2(N656), .ZN(n567) );
  nd12d0 U568 ( .A1(n573), .A2(n572), .ZN(N852) );
  nd12d0 U569 ( .A1(n571), .A2(n570), .ZN(n573) );
  nd12d0 U570 ( .A1(n6), .A2(N657), .ZN(n572) );
  nd12d0 U571 ( .A1(n578), .A2(n577), .ZN(N853) );
  nd12d0 U572 ( .A1(n576), .A2(n575), .ZN(n578) );
  nd12d0 U573 ( .A1(n6), .A2(N658), .ZN(n577) );
  nd12d0 U574 ( .A1(n583), .A2(n582), .ZN(N854) );
  nd12d0 U575 ( .A1(n581), .A2(n580), .ZN(n583) );
  nd12d0 U576 ( .A1(n7), .A2(N659), .ZN(n582) );
  nd12d0 U577 ( .A1(n588), .A2(n587), .ZN(N855) );
  nd12d0 U578 ( .A1(n586), .A2(n585), .ZN(n588) );
  nd12d0 U579 ( .A1(n7), .A2(N660), .ZN(n587) );
  nd12d0 U580 ( .A1(n593), .A2(n592), .ZN(N856) );
  nd12d0 U581 ( .A1(n591), .A2(n590), .ZN(n593) );
  nd12d0 U582 ( .A1(n7), .A2(N661), .ZN(n592) );
  nd12d0 U583 ( .A1(n598), .A2(n597), .ZN(N857) );
  nd12d0 U584 ( .A1(n596), .A2(n595), .ZN(n598) );
  nd12d0 U585 ( .A1(n7), .A2(N662), .ZN(n597) );
  nd12d0 U586 ( .A1(n603), .A2(n602), .ZN(N858) );
  nd12d0 U587 ( .A1(n601), .A2(n600), .ZN(n603) );
  nd12d0 U588 ( .A1(n6), .A2(N663), .ZN(n602) );
  nd12d0 U589 ( .A1(n613), .A2(n612), .ZN(N860) );
  nd12d0 U590 ( .A1(n611), .A2(n610), .ZN(n613) );
  nd12d0 U591 ( .A1(n6), .A2(N665), .ZN(n612) );
  nd12d0 U592 ( .A1(n703), .A2(n702), .ZN(N888) );
  nd12d0 U593 ( .A1(n701), .A2(n700), .ZN(n703) );
  nd12d0 U594 ( .A1(n7), .A2(N725), .ZN(n702) );
  nd12d0 U595 ( .A1(n708), .A2(n707), .ZN(N889) );
  nd12d0 U596 ( .A1(n706), .A2(n705), .ZN(n708) );
  nd12d0 U597 ( .A1(n7), .A2(N726), .ZN(n707) );
  nd12d0 U598 ( .A1(n538), .A2(n537), .ZN(N845) );
  nd12d0 U599 ( .A1(n536), .A2(n535), .ZN(n538) );
  nd12d0 U600 ( .A1(n7), .A2(N650), .ZN(n537) );
  nd12d0 U601 ( .A1(n543), .A2(n542), .ZN(N846) );
  nd12d0 U602 ( .A1(n541), .A2(n540), .ZN(n543) );
  nd12d0 U603 ( .A1(n6), .A2(N651), .ZN(n542) );
  nd12d0 U604 ( .A1(n548), .A2(n547), .ZN(N847) );
  nd12d0 U605 ( .A1(n546), .A2(n545), .ZN(n548) );
  nd12d0 U606 ( .A1(n7), .A2(N652), .ZN(n547) );
  nd12d0 U607 ( .A1(n553), .A2(n552), .ZN(N848) );
  nd12d0 U608 ( .A1(n551), .A2(n550), .ZN(n553) );
  nd12d0 U609 ( .A1(n6), .A2(N653), .ZN(n552) );
  nd12d0 U610 ( .A1(n558), .A2(n557), .ZN(N849) );
  nd12d0 U611 ( .A1(n556), .A2(n555), .ZN(n558) );
  nd12d0 U612 ( .A1(n7), .A2(N654), .ZN(n557) );
  nd12d0 U613 ( .A1(n643), .A2(n642), .ZN(N876) );
  nd12d0 U614 ( .A1(n641), .A2(n640), .ZN(n643) );
  nd12d0 U615 ( .A1(n7), .A2(N713), .ZN(n642) );
  nd12d0 U616 ( .A1(n648), .A2(n647), .ZN(N877) );
  nd12d0 U617 ( .A1(n646), .A2(n645), .ZN(n648) );
  nd12d0 U618 ( .A1(n6), .A2(N714), .ZN(n647) );
  nd12d0 U619 ( .A1(n653), .A2(n652), .ZN(N878) );
  nd12d0 U620 ( .A1(n651), .A2(n650), .ZN(n653) );
  nd12d0 U621 ( .A1(n7), .A2(N715), .ZN(n652) );
  nd12d0 U622 ( .A1(n658), .A2(n657), .ZN(N879) );
  nd12d0 U623 ( .A1(n656), .A2(n655), .ZN(n658) );
  nd12d0 U624 ( .A1(n6), .A2(N716), .ZN(n657) );
  nd12d0 U625 ( .A1(n663), .A2(n662), .ZN(N880) );
  nd12d0 U626 ( .A1(n661), .A2(n660), .ZN(n663) );
  nd12d0 U627 ( .A1(n6), .A2(N717), .ZN(n662) );
  nd12d0 U628 ( .A1(n668), .A2(n667), .ZN(N881) );
  nd12d0 U629 ( .A1(n666), .A2(n665), .ZN(n668) );
  nd12d0 U630 ( .A1(n6), .A2(N718), .ZN(n667) );
  nd12d0 U631 ( .A1(n523), .A2(n522), .ZN(N842) );
  nd12d0 U632 ( .A1(n521), .A2(n520), .ZN(n523) );
  nd12d0 U633 ( .A1(n6), .A2(N647), .ZN(n522) );
  nd12d0 U634 ( .A1(n528), .A2(n527), .ZN(N843) );
  nd12d0 U635 ( .A1(n526), .A2(n525), .ZN(n528) );
  nd12d0 U693 ( .A1(n7), .A2(N648), .ZN(n527) );
  nd12d0 U702 ( .A1(n533), .A2(n532), .ZN(N844) );
  nd12d0 U703 ( .A1(n531), .A2(n530), .ZN(n533) );
  nd12d0 U753 ( .A1(n6), .A2(N649), .ZN(n532) );
  nd12d0 U756 ( .A1(n633), .A2(n632), .ZN(N874) );
  nd12d0 U757 ( .A1(n631), .A2(n630), .ZN(n633) );
  nd12d0 U758 ( .A1(n7), .A2(N711), .ZN(n632) );
  nd12d0 U759 ( .A1(n638), .A2(n637), .ZN(N875) );
  nd12d0 U760 ( .A1(n636), .A2(n635), .ZN(n638) );
  nd12d0 U761 ( .A1(n6), .A2(N712), .ZN(n637) );
  nd12d0 U762 ( .A1(n519), .A2(n5), .ZN(n13) );
  nd12d0 U763 ( .A1(n519), .A2(n5), .ZN(n14) );
  nd12d0 U764 ( .A1(n519), .A2(n5), .ZN(n736) );
  an12d1 U765 ( .A2(n484), .A1(n492), .Z(n499) );
  an12d1 U766 ( .A2(n484), .A1(n493), .Z(n500) );
  an12d1 U767 ( .A2(n484), .A1(n493), .Z(n479) );
  nr02d0 U768 ( .A1(n494), .A2(n484), .ZN(n478) );
  nr02d0 U769 ( .A1(n492), .A2(n484), .ZN(n497) );
  nr02d0 U770 ( .A1(n494), .A2(n484), .ZN(n498) );
  an02d1 U771 ( .A1(n5), .A2(n519), .Z(n1) );
  bufbd1 U772 ( .I(n942), .Z(n16) );
  bufbd1 U773 ( .I(n942), .Z(n15) );
  inv0d1 U774 ( .I(n474), .ZN(n483) );
  nd12d0 U775 ( .A1(n740), .A2(n16), .ZN(n474) );
  an02d1 U776 ( .A1(n492), .A2(n946), .Z(n2) );
  bufbd1 U777 ( .I(n467), .Z(n508) );
  bufbd1 U778 ( .I(n467), .Z(n509) );
  bufbd1 U779 ( .I(n467), .Z(n510) );
  bufbd1 U780 ( .I(n467), .Z(n511) );
  bufbd1 U781 ( .I(n467), .Z(n512) );
  bufbd1 U782 ( .I(n467), .Z(n513) );
  an02d1 U783 ( .A1(n15), .A2(n740), .Z(n3) );
  an02d1 U784 ( .A1(n15), .A2(n740), .Z(n4) );
  nd12d0 U785 ( .A1(n13), .A2(N738), .ZN(n520) );
  bufbd1 U786 ( .I(n467), .Z(n514) );
  nd12d0 U787 ( .A1(n13), .A2(N762), .ZN(n630) );
  nd12d0 U788 ( .A1(n765), .A2(n764), .ZN(N545) );
  nd12d0 U789 ( .A1(n16), .A2(N350), .ZN(n764) );
  nd12d0 U790 ( .A1(n763), .A2(n762), .ZN(n765) );
  nd12d0 U791 ( .A1(n760), .A2(n759), .ZN(N544) );
  nd12d0 U792 ( .A1(n15), .A2(N349), .ZN(n759) );
  nd12d0 U793 ( .A1(n758), .A2(n757), .ZN(n760) );
  nd12d0 U794 ( .A1(n490), .A2(N416), .ZN(n757) );
  inv0d1 U795 ( .I(n491), .ZN(n492) );
  inv0d1 U796 ( .I(n491), .ZN(n493) );
  inv0d1 U797 ( .I(n491), .ZN(n494) );
  nd12d0 U798 ( .A1(n9), .A2(s3_op2[27]), .ZN(n726) );
  nd12d0 U799 ( .A1(n14), .A2(N781), .ZN(n725) );
  nd12d0 U800 ( .A1(n6), .A2(N730), .ZN(n724) );
  nd12d0 U801 ( .A1(n10), .A2(s3_op2[28]), .ZN(n729) );
  nd12d0 U802 ( .A1(n736), .A2(N782), .ZN(n728) );
  nd12d0 U803 ( .A1(n5), .A2(N731), .ZN(n727) );
  nd12d0 U804 ( .A1(n10), .A2(s3_op2[29]), .ZN(n732) );
  nd12d0 U805 ( .A1(n13), .A2(N783), .ZN(n731) );
  nd12d0 U806 ( .A1(n7), .A2(N732), .ZN(n730) );
  nd12d0 U807 ( .A1(n11), .A2(s3_op2[30]), .ZN(n735) );
  nd12d0 U808 ( .A1(n14), .A2(N784), .ZN(n734) );
  nd12d0 U809 ( .A1(n6), .A2(N733), .ZN(n733) );
  nd12d0 U810 ( .A1(n12), .A2(s3_op2[31]), .ZN(n739) );
  nd12d0 U811 ( .A1(n736), .A2(N785), .ZN(n738) );
  nd02d1 U812 ( .A1(N734), .A2(n2), .ZN(n737) );
  nd12d0 U813 ( .A1(n12), .A2(s3_op1[27]), .ZN(n616) );
  nd12d0 U814 ( .A1(n14), .A2(N757), .ZN(n615) );
  nd12d0 U815 ( .A1(n7), .A2(N666), .ZN(n614) );
  nd12d0 U816 ( .A1(n8), .A2(s3_op1[28]), .ZN(n619) );
  nd12d0 U817 ( .A1(n736), .A2(N758), .ZN(n618) );
  nd12d0 U818 ( .A1(n6), .A2(N667), .ZN(n617) );
  nd12d0 U819 ( .A1(n12), .A2(s3_op1[29]), .ZN(n622) );
  nd12d0 U820 ( .A1(n13), .A2(N759), .ZN(n621) );
  nd12d0 U821 ( .A1(n7), .A2(N668), .ZN(n620) );
  nd12d0 U822 ( .A1(n8), .A2(s3_op1[30]), .ZN(n625) );
  nd12d0 U823 ( .A1(n14), .A2(N760), .ZN(n624) );
  nd12d0 U824 ( .A1(n6), .A2(N669), .ZN(n623) );
  nd12d0 U825 ( .A1(n9), .A2(s3_op1[31]), .ZN(n628) );
  nd12d0 U826 ( .A1(n736), .A2(N761), .ZN(n627) );
  nd02d1 U827 ( .A1(N670), .A2(n2), .ZN(n626) );
  nd12d0 U828 ( .A1(n471), .A2(s2_op1[31]), .ZN(n846) );
  nd12d0 U829 ( .A1(n15), .A2(N377), .ZN(n844) );
  nd12d0 U830 ( .A1(n475), .A2(N444), .ZN(n845) );
  nd12d0 U831 ( .A1(n473), .A2(s2_op2[29]), .ZN(n938) );
  nd12d0 U832 ( .A1(n476), .A2(N474), .ZN(n937) );
  nd12d0 U833 ( .A1(n15), .A2(N407), .ZN(n936) );
  nd12d0 U834 ( .A1(n17), .A2(s2_op2[30]), .ZN(n941) );
  nd12d0 U835 ( .A1(n477), .A2(N475), .ZN(n940) );
  nd12d0 U836 ( .A1(n942), .A2(N408), .ZN(n939) );
  nd12d0 U837 ( .A1(n473), .A2(s2_op1[25]), .ZN(n828) );
  nd12d0 U838 ( .A1(n16), .A2(N371), .ZN(n826) );
  nd12d0 U839 ( .A1(n488), .A2(N438), .ZN(n827) );
  nd12d0 U840 ( .A1(n17), .A2(s2_op1[26]), .ZN(n831) );
  nd12d0 U841 ( .A1(n942), .A2(N372), .ZN(n829) );
  nd12d0 U842 ( .A1(n477), .A2(N439), .ZN(n830) );
  nd12d0 U843 ( .A1(n468), .A2(s2_op1[27]), .ZN(n834) );
  nd12d0 U844 ( .A1(n15), .A2(N373), .ZN(n832) );
  nd12d0 U845 ( .A1(n486), .A2(N440), .ZN(n833) );
  nd12d0 U846 ( .A1(n472), .A2(s2_op1[28]), .ZN(n837) );
  nd12d0 U847 ( .A1(n16), .A2(N374), .ZN(n835) );
  nd12d0 U848 ( .A1(n489), .A2(N441), .ZN(n836) );
  nd12d0 U849 ( .A1(n473), .A2(s2_op1[29]), .ZN(n840) );
  nd12d0 U850 ( .A1(n15), .A2(N375), .ZN(n838) );
  nd12d0 U851 ( .A1(n489), .A2(N442), .ZN(n839) );
  nd12d0 U852 ( .A1(n470), .A2(s2_op1[30]), .ZN(n843) );
  nd12d0 U853 ( .A1(n16), .A2(N376), .ZN(n841) );
  nd12d0 U854 ( .A1(n490), .A2(N443), .ZN(n842) );
  nd12d0 U855 ( .A1(n468), .A2(s2_op2[31]), .ZN(n945) );
  nd12d0 U856 ( .A1(n485), .A2(N476), .ZN(n944) );
  nd12d0 U857 ( .A1(n16), .A2(N409), .ZN(n943) );
  nd12d0 U858 ( .A1(n17), .A2(s2_op2[22]), .ZN(n917) );
  nd12d0 U859 ( .A1(n488), .A2(N467), .ZN(n916) );
  nd12d0 U860 ( .A1(n16), .A2(N400), .ZN(n915) );
  nd12d0 U861 ( .A1(n470), .A2(s2_op2[24]), .ZN(n923) );
  nd12d0 U862 ( .A1(n489), .A2(N469), .ZN(n922) );
  nd12d0 U863 ( .A1(n16), .A2(N402), .ZN(n921) );
  nd12d0 U864 ( .A1(n471), .A2(s2_op2[25]), .ZN(n926) );
  nd12d0 U865 ( .A1(n476), .A2(N470), .ZN(n925) );
  nd12d0 U866 ( .A1(n15), .A2(N403), .ZN(n924) );
  nd12d0 U867 ( .A1(n470), .A2(s2_op2[26]), .ZN(n929) );
  nd12d0 U868 ( .A1(n489), .A2(N471), .ZN(n928) );
  nd12d0 U869 ( .A1(n16), .A2(N404), .ZN(n927) );
  nd12d0 U870 ( .A1(n471), .A2(s2_op2[27]), .ZN(n932) );
  nd12d0 U871 ( .A1(n490), .A2(N472), .ZN(n931) );
  nd12d0 U872 ( .A1(n942), .A2(N405), .ZN(n930) );
  nd12d0 U873 ( .A1(n472), .A2(s2_op2[28]), .ZN(n935) );
  nd12d0 U874 ( .A1(n475), .A2(N473), .ZN(n934) );
  nd12d0 U875 ( .A1(n15), .A2(N406), .ZN(n933) );
  nd12d0 U876 ( .A1(n471), .A2(s2_op1[23]), .ZN(n822) );
  nd12d0 U877 ( .A1(n942), .A2(N369), .ZN(n820) );
  nd12d0 U878 ( .A1(n486), .A2(N436), .ZN(n821) );
  nd12d0 U879 ( .A1(n472), .A2(s2_op1[24]), .ZN(n825) );
  nd12d0 U880 ( .A1(n15), .A2(N370), .ZN(n823) );
  nd12d0 U881 ( .A1(n487), .A2(N437), .ZN(n824) );
  mx02d0 U882 ( .I0(s3_op1[6]), .I1(N645), .S(n2), .Z(N840) );
  mx02d0 U883 ( .I0(s3_op1[7]), .I1(N646), .S(n2), .Z(N841) );
  mx02d0 U884 ( .I0(s3_op2[6]), .I1(N709), .S(n2), .Z(N872) );
  mx02d0 U885 ( .I0(s3_op2[7]), .I1(N710), .S(n2), .Z(N873) );
  nd12d0 U886 ( .A1(n470), .A2(s2_op1[20]), .ZN(n813) );
  nd12d0 U887 ( .A1(n942), .A2(N366), .ZN(n811) );
  nd12d0 U888 ( .A1(n476), .A2(N433), .ZN(n812) );
  nd12d0 U889 ( .A1(n471), .A2(s2_op1[21]), .ZN(n816) );
  nd12d0 U890 ( .A1(n15), .A2(N367), .ZN(n814) );
  nd12d0 U891 ( .A1(n477), .A2(N434), .ZN(n815) );
  nd12d0 U892 ( .A1(n470), .A2(s2_op1[22]), .ZN(n819) );
  nd12d0 U893 ( .A1(n16), .A2(N368), .ZN(n817) );
  nd12d0 U894 ( .A1(n485), .A2(N435), .ZN(n818) );
  nd12d0 U895 ( .A1(n468), .A2(s2_op2[23]), .ZN(n920) );
  nd12d0 U896 ( .A1(n487), .A2(N468), .ZN(n919) );
  nd12d0 U897 ( .A1(n942), .A2(N401), .ZN(n918) );
  nd12d0 U898 ( .A1(n471), .A2(s2_op2[17]), .ZN(n902) );
  nd12d0 U899 ( .A1(n476), .A2(N462), .ZN(n901) );
  nd12d0 U900 ( .A1(n15), .A2(N395), .ZN(n900) );
  nd12d0 U901 ( .A1(n472), .A2(s2_op2[18]), .ZN(n905) );
  nd12d0 U902 ( .A1(n477), .A2(N463), .ZN(n904) );
  nd12d0 U903 ( .A1(n16), .A2(N396), .ZN(n903) );
  nd12d0 U904 ( .A1(n17), .A2(s2_op2[20]), .ZN(n911) );
  nd12d0 U905 ( .A1(n486), .A2(N465), .ZN(n910) );
  nd12d0 U906 ( .A1(n15), .A2(N398), .ZN(n909) );
  nd12d0 U907 ( .A1(n473), .A2(s2_op1[15]), .ZN(n798) );
  nd12d0 U908 ( .A1(n15), .A2(N361), .ZN(n796) );
  nd12d0 U909 ( .A1(n490), .A2(N428), .ZN(n797) );
  nd12d0 U910 ( .A1(n17), .A2(s2_op1[16]), .ZN(n801) );
  nd12d0 U911 ( .A1(n16), .A2(N362), .ZN(n799) );
  nd12d0 U912 ( .A1(n475), .A2(N429), .ZN(n800) );
  nd12d0 U913 ( .A1(n468), .A2(s2_op1[19]), .ZN(n810) );
  nd12d0 U914 ( .A1(n16), .A2(N365), .ZN(n808) );
  nd12d0 U915 ( .A1(n488), .A2(N432), .ZN(n809) );
  mx02d0 U916 ( .I0(s3_op1[3]), .I1(N642), .S(n2), .Z(N837) );
  mx02d0 U917 ( .I0(s3_op1[4]), .I1(N643), .S(n2), .Z(N838) );
  mx02d0 U918 ( .I0(s3_op1[5]), .I1(N644), .S(n2), .Z(N839) );
  mx02d0 U919 ( .I0(s3_op2[3]), .I1(N706), .S(n2), .Z(N869) );
  mx02d0 U920 ( .I0(s3_op2[4]), .I1(N707), .S(n2), .Z(N870) );
  mx02d0 U921 ( .I0(s3_op2[5]), .I1(N708), .S(n2), .Z(N871) );
  nd12d0 U922 ( .A1(n468), .A2(s2_op1[17]), .ZN(n804) );
  nd12d0 U923 ( .A1(n942), .A2(N363), .ZN(n802) );
  nd12d0 U924 ( .A1(n476), .A2(N430), .ZN(n803) );
  nd12d0 U925 ( .A1(n17), .A2(s2_op1[18]), .ZN(n807) );
  nd12d0 U926 ( .A1(n15), .A2(N364), .ZN(n805) );
  nd12d0 U927 ( .A1(n485), .A2(N431), .ZN(n806) );
  nd12d0 U928 ( .A1(n470), .A2(s2_op2[16]), .ZN(n899) );
  nd12d0 U929 ( .A1(n475), .A2(N461), .ZN(n898) );
  nd12d0 U930 ( .A1(n942), .A2(N394), .ZN(n897) );
  nd12d0 U931 ( .A1(n473), .A2(s2_op2[19]), .ZN(n908) );
  nd12d0 U932 ( .A1(n485), .A2(N464), .ZN(n907) );
  nd12d0 U933 ( .A1(n942), .A2(N397), .ZN(n906) );
  nd12d0 U934 ( .A1(n468), .A2(s2_op2[21]), .ZN(n914) );
  nd12d0 U935 ( .A1(n487), .A2(N466), .ZN(n913) );
  nd12d0 U936 ( .A1(n942), .A2(N399), .ZN(n912) );
  nd12d0 U937 ( .A1(n473), .A2(s2_op2[11]), .ZN(n884) );
  nd12d0 U938 ( .A1(n489), .A2(N456), .ZN(n883) );
  nd12d0 U939 ( .A1(n15), .A2(N389), .ZN(n882) );
  nd12d0 U940 ( .A1(n17), .A2(s2_op2[12]), .ZN(n887) );
  nd12d0 U941 ( .A1(n490), .A2(N457), .ZN(n886) );
  nd12d0 U942 ( .A1(n16), .A2(N390), .ZN(n885) );
  nd12d0 U943 ( .A1(n468), .A2(s2_op2[13]), .ZN(n890) );
  nd12d0 U944 ( .A1(n475), .A2(N458), .ZN(n889) );
  nd12d0 U945 ( .A1(n16), .A2(N391), .ZN(n888) );
  nd12d0 U946 ( .A1(n472), .A2(s2_op2[14]), .ZN(n893) );
  nd12d0 U947 ( .A1(n486), .A2(N459), .ZN(n892) );
  nd12d0 U948 ( .A1(n15), .A2(N392), .ZN(n891) );
  nd12d0 U949 ( .A1(n471), .A2(s2_op2[9]), .ZN(n878) );
  nd12d0 U950 ( .A1(n487), .A2(N454), .ZN(n877) );
  nd12d0 U951 ( .A1(n16), .A2(N387), .ZN(n876) );
  nd12d0 U952 ( .A1(n472), .A2(s2_op1[10]), .ZN(n783) );
  nd12d0 U953 ( .A1(n16), .A2(N356), .ZN(n781) );
  nd12d0 U954 ( .A1(n487), .A2(N423), .ZN(n782) );
  nd12d0 U955 ( .A1(n468), .A2(s2_op1[9]), .ZN(n780) );
  nd12d0 U956 ( .A1(n15), .A2(N355), .ZN(n778) );
  nd12d0 U957 ( .A1(n477), .A2(N422), .ZN(n779) );
  nd12d0 U958 ( .A1(n473), .A2(s2_op1[11]), .ZN(n786) );
  nd12d0 U959 ( .A1(n942), .A2(N357), .ZN(n784) );
  nd12d0 U960 ( .A1(n486), .A2(N424), .ZN(n785) );
  nd12d0 U961 ( .A1(n470), .A2(s2_op1[12]), .ZN(n789) );
  nd12d0 U962 ( .A1(n15), .A2(N358), .ZN(n787) );
  nd12d0 U963 ( .A1(n487), .A2(N425), .ZN(n788) );
  mx02d0 U964 ( .I0(s3_op1[1]), .I1(N640), .S(n2), .Z(N835) );
  mx02d0 U965 ( .I0(s3_op1[2]), .I1(N641), .S(n2), .Z(N836) );
  mx02d0 U966 ( .I0(s3_op2[1]), .I1(N704), .S(n2), .Z(N867) );
  mx02d0 U967 ( .I0(s3_op2[2]), .I1(N705), .S(n2), .Z(N868) );
  nd12d0 U968 ( .A1(n471), .A2(s2_op1[13]), .ZN(n792) );
  nd12d0 U969 ( .A1(n16), .A2(N359), .ZN(n790) );
  nd12d0 U970 ( .A1(n488), .A2(N426), .ZN(n791) );
  nd12d0 U971 ( .A1(n472), .A2(s2_op1[14]), .ZN(n795) );
  nd12d0 U972 ( .A1(n942), .A2(N360), .ZN(n793) );
  nd12d0 U973 ( .A1(n489), .A2(N427), .ZN(n794) );
  nd12d0 U974 ( .A1(n471), .A2(s2_op2[7]), .ZN(n872) );
  nd12d0 U975 ( .A1(n490), .A2(N452), .ZN(n871) );
  nd12d0 U976 ( .A1(n942), .A2(N385), .ZN(n870) );
  nd12d0 U977 ( .A1(n472), .A2(s2_op2[10]), .ZN(n881) );
  nd12d0 U978 ( .A1(n488), .A2(N455), .ZN(n880) );
  nd12d0 U979 ( .A1(n942), .A2(N388), .ZN(n879) );
  nd12d0 U980 ( .A1(n473), .A2(s2_op2[15]), .ZN(n896) );
  nd12d0 U981 ( .A1(n488), .A2(N460), .ZN(n895) );
  nd12d0 U982 ( .A1(n942), .A2(N393), .ZN(n894) );
  nd12d0 U983 ( .A1(n517), .A2(trans2), .ZN(n467) );
  nr02d0 U984 ( .A1(n440), .A2(n494), .ZN(n482) );
  nd02d1 U985 ( .A1(n515), .A2(trans2), .ZN(n740) );
  nd12d0 U986 ( .A1(n470), .A2(s2_op2[6]), .ZN(n869) );
  nd12d0 U987 ( .A1(n487), .A2(N451), .ZN(n868) );
  nd12d0 U988 ( .A1(n16), .A2(N384), .ZN(n867) );
  nd12d0 U989 ( .A1(n472), .A2(s2_op1[6]), .ZN(n771) );
  nd12d0 U990 ( .A1(n477), .A2(N419), .ZN(n770) );
  nd12d0 U991 ( .A1(n15), .A2(N352), .ZN(n769) );
  nd12d0 U992 ( .A1(n17), .A2(s2_op2[4]), .ZN(n863) );
  nd12d0 U993 ( .A1(n485), .A2(N449), .ZN(n862) );
  nd12d0 U994 ( .A1(n942), .A2(N382), .ZN(n861) );
  nd12d0 U995 ( .A1(n473), .A2(s2_op1[7]), .ZN(n774) );
  nd12d0 U996 ( .A1(n485), .A2(N420), .ZN(n773) );
  nd12d0 U997 ( .A1(n16), .A2(N353), .ZN(n772) );
  nd12d0 U998 ( .A1(n468), .A2(s2_op2[5]), .ZN(n866) );
  nd12d0 U999 ( .A1(n485), .A2(N450), .ZN(n865) );
  nd12d0 U1000 ( .A1(n15), .A2(N383), .ZN(n864) );
  nd12d0 U1001 ( .A1(n16), .A2(N381), .ZN(n858) );
  nd12d0 U1002 ( .A1(n468), .A2(s2_op2[3]), .ZN(n860) );
  nd12d0 U1003 ( .A1(n477), .A2(N448), .ZN(n859) );
  nd12d0 U1004 ( .A1(n15), .A2(N380), .ZN(n855) );
  nd12d0 U1005 ( .A1(n17), .A2(s2_op2[2]), .ZN(n857) );
  nd12d0 U1006 ( .A1(n476), .A2(N447), .ZN(n856) );
  nd12d0 U1007 ( .A1(n471), .A2(s2_op1[5]), .ZN(n768) );
  nd12d0 U1008 ( .A1(n476), .A2(N418), .ZN(n767) );
  nd12d0 U1009 ( .A1(n942), .A2(N351), .ZN(n766) );
  nd12d0 U1010 ( .A1(n470), .A2(s2_op2[8]), .ZN(n875) );
  nd12d0 U1011 ( .A1(n486), .A2(N453), .ZN(n874) );
  nd12d0 U1012 ( .A1(n15), .A2(N386), .ZN(n873) );
  nd12d0 U1013 ( .A1(n17), .A2(s2_op1[8]), .ZN(n777) );
  nd12d0 U1014 ( .A1(n942), .A2(N354), .ZN(n775) );
  nd12d0 U1015 ( .A1(n475), .A2(N421), .ZN(n776) );
  nr02d0 U1016 ( .A1(n517), .A2(trans2), .ZN(n495) );
  nr02d0 U1017 ( .A1(n517), .A2(trans2), .ZN(n496) );
  nd02d1 U1018 ( .A1(trans2), .A2(trans3), .ZN(n519) );
  nr02d0 U1019 ( .A1(n517), .A2(trans2), .ZN(n469) );
  inv0d1 U1020 ( .I(operation[2]), .ZN(n460) );
  inv0d1 U1021 ( .I(operation[3]), .ZN(n464) );
  bufbd1 U1022 ( .I(trans1), .Z(n516) );
  inv0d1 U1023 ( .I(operation[1]), .ZN(n463) );
  bufbd1 U1024 ( .I(n480), .Z(n501) );
  bufbd1 U1025 ( .I(trans1), .Z(n515) );
  inv0d1 U1026 ( .I(operation[0]), .ZN(n466) );
  nd12d0 U1027 ( .A1(n461), .A2(n462), .ZN(c_trans1) );
  inv0d1 U1028 ( .I(rem_red), .ZN(n491) );
  xr03d1 U1029 ( .A1(s4_op1[1]), .A2(s4_op1[0]), .A3(n458), .Z(s5_result[0])
         );
  xr03d1 U1030 ( .A1(s4_op1[3]), .A2(s4_op1[2]), .A3(n451), .Z(s5_result[1])
         );
  xr03d1 U1031 ( .A1(s4_op1[5]), .A2(s4_op1[4]), .A3(n450), .Z(s5_result[2])
         );
  xr03d1 U1032 ( .A1(s4_op1[7]), .A2(s4_op1[6]), .A3(n449), .Z(s5_result[3])
         );
  xr03d1 U1033 ( .A1(s4_op1[9]), .A2(s4_op1[8]), .A3(n448), .Z(s5_result[4])
         );
  xr03d1 U1034 ( .A1(s4_op1[11]), .A2(s4_op1[10]), .A3(n447), .Z(s5_result[5])
         );
  xr03d1 U1035 ( .A1(s4_op1[13]), .A2(s4_op1[12]), .A3(n446), .Z(s5_result[6])
         );
  xr03d1 U1036 ( .A1(s4_op1[15]), .A2(s4_op1[14]), .A3(n445), .Z(s5_result[7])
         );
  xr03d1 U1037 ( .A1(s4_op1[17]), .A2(s4_op1[16]), .A3(n444), .Z(s5_result[8])
         );
  xr03d1 U1038 ( .A1(s4_op1[19]), .A2(s4_op1[18]), .A3(n443), .Z(s5_result[9])
         );
  xr03d1 U1039 ( .A1(s4_op1[21]), .A2(s4_op1[20]), .A3(n457), .Z(s5_result[10]) );
  xr03d1 U1040 ( .A1(s4_op1[23]), .A2(s4_op1[22]), .A3(n456), .Z(s5_result[11]) );
  xr03d1 U1041 ( .A1(s4_op1[25]), .A2(s4_op1[24]), .A3(n455), .Z(s5_result[12]) );
  xr03d1 U1042 ( .A1(s4_op1[27]), .A2(s4_op1[26]), .A3(n454), .Z(s5_result[13]) );
  xr03d1 U1043 ( .A1(s4_op1[29]), .A2(s4_op1[28]), .A3(n453), .Z(s5_result[14]) );
  xr03d1 U1044 ( .A1(s4_op1[31]), .A2(s4_op1[30]), .A3(n452), .Z(s5_result[15]) );
  nd12d0 U1045 ( .A1(n475), .A2(N417), .ZN(n762) );
  nd12d0 U1046 ( .A1(n755), .A2(n754), .ZN(N543) );
  nd12d0 U1047 ( .A1(n942), .A2(N348), .ZN(n754) );
  nd12d0 U1048 ( .A1(n753), .A2(n752), .ZN(n755) );
  nd12d0 U1049 ( .A1(n489), .A2(N415), .ZN(n752) );
  nd12d0 U1050 ( .A1(n16), .A2(N347), .ZN(n750) );
  bufbd1 U1051 ( .I(trans1), .Z(n517) );
  nd12d0 U1052 ( .A1(n470), .A2(s2_op1[0]), .ZN(n744) );
  nd12d0 U1053 ( .A1(n741), .A2(n851), .ZN(n743) );
  nd12d0 U1054 ( .A1(n472), .A2(s2_op2[0]), .ZN(n850) );
  nd12d0 U1055 ( .A1(n847), .A2(n851), .ZN(n849) );
  mx02d0 U1056 ( .I0(s3_op1[0]), .I1(N639), .S(n2), .Z(N834) );
  mx02d0 U1057 ( .I0(s3_op2[0]), .I1(N703), .S(n2), .Z(N866) );
  nd12d0 U1058 ( .A1(n942), .A2(N379), .ZN(n852) );
  nd12d0 U1059 ( .A1(n473), .A2(s2_op2[1]), .ZN(n854) );
  inv0d1 U1060 ( .I(s3_op2[16]), .ZN(n669) );
  inv0d1 U1061 ( .I(s3_op1[11]), .ZN(n534) );
  inv0d1 U1062 ( .I(s3_op1[12]), .ZN(n539) );
  inv0d1 U1063 ( .I(s3_op1[13]), .ZN(n544) );
  inv0d1 U1064 ( .I(s3_op1[14]), .ZN(n549) );
  inv0d1 U1065 ( .I(trans3), .ZN(n942) );
  inv0d1 U1066 ( .I(s3_op1[8]), .ZN(n518) );
  inv0d1 U1067 ( .I(s3_op1[9]), .ZN(n524) );
  inv0d1 U1068 ( .I(s3_op1[15]), .ZN(n554) );
  inv0d1 U1069 ( .I(s3_op2[8]), .ZN(n629) );
  inv0d1 U1070 ( .I(s3_op2[9]), .ZN(n634) );
  inv0d1 U1071 ( .I(s3_op2[11]), .ZN(n644) );
  inv0d1 U1072 ( .I(s3_op2[12]), .ZN(n649) );
  inv0d1 U1073 ( .I(s3_op2[13]), .ZN(n654) );
  inv0d1 U1074 ( .I(s3_op2[14]), .ZN(n659) );
  inv0d1 U1075 ( .I(s3_op2[15]), .ZN(n664) );
  inv0d1 U1076 ( .I(s3_op1[10]), .ZN(n529) );
  inv0d1 U1077 ( .I(s3_op2[10]), .ZN(n639) );
  inv0d1 U1078 ( .I(n440), .ZN(n946) );
  nr02d0 U1079 ( .A1(n8), .A2(n518), .ZN(n521) );
  nr02d0 U1080 ( .A1(n9), .A2(n524), .ZN(n526) );
  nr02d0 U1081 ( .A1(n10), .A2(n529), .ZN(n531) );
  nr02d0 U1082 ( .A1(n8), .A2(n534), .ZN(n536) );
  nr02d0 U1083 ( .A1(n9), .A2(n539), .ZN(n541) );
  nr02d0 U1084 ( .A1(n11), .A2(n544), .ZN(n546) );
  nr02d0 U1085 ( .A1(n12), .A2(n549), .ZN(n551) );
  nr02d0 U1086 ( .A1(n8), .A2(n554), .ZN(n556) );
  inv0d1 U1087 ( .I(s3_op1[16]), .ZN(n559) );
  nr02d0 U1088 ( .A1(n10), .A2(n559), .ZN(n561) );
  inv0d1 U1089 ( .I(s3_op1[17]), .ZN(n564) );
  nr02d0 U1090 ( .A1(n11), .A2(n564), .ZN(n566) );
  inv0d1 U1091 ( .I(s3_op1[18]), .ZN(n569) );
  nr02d0 U1092 ( .A1(n9), .A2(n569), .ZN(n571) );
  inv0d1 U1093 ( .I(s3_op1[19]), .ZN(n574) );
  nr02d0 U1094 ( .A1(n10), .A2(n574), .ZN(n576) );
  inv0d1 U1095 ( .I(s3_op1[20]), .ZN(n579) );
  nr02d0 U1096 ( .A1(n11), .A2(n579), .ZN(n581) );
  inv0d1 U1097 ( .I(s3_op1[21]), .ZN(n584) );
  nr02d0 U1098 ( .A1(n12), .A2(n584), .ZN(n586) );
  inv0d1 U1099 ( .I(s3_op1[22]), .ZN(n589) );
  nr02d0 U1100 ( .A1(n8), .A2(n589), .ZN(n591) );
  inv0d1 U1101 ( .I(s3_op1[23]), .ZN(n594) );
  nr02d0 U1102 ( .A1(n12), .A2(n594), .ZN(n596) );
  inv0d1 U1103 ( .I(s3_op1[24]), .ZN(n599) );
  nr02d0 U1104 ( .A1(n8), .A2(n599), .ZN(n601) );
  inv0d1 U1105 ( .I(s3_op1[25]), .ZN(n604) );
  nr02d0 U1106 ( .A1(n9), .A2(n604), .ZN(n606) );
  inv0d1 U1107 ( .I(s3_op1[26]), .ZN(n609) );
  nr02d0 U1108 ( .A1(n9), .A2(n609), .ZN(n611) );
  nd03d0 U1109 ( .A1(n616), .A2(n615), .A3(n614), .ZN(N861) );
  nd03d0 U1110 ( .A1(n619), .A2(n618), .A3(n617), .ZN(N862) );
  nd03d0 U1111 ( .A1(n622), .A2(n621), .A3(n620), .ZN(N863) );
  nd03d0 U1112 ( .A1(n625), .A2(n624), .A3(n623), .ZN(N864) );
  nd03d0 U1113 ( .A1(n628), .A2(n627), .A3(n626), .ZN(N865) );
  nr02d0 U1114 ( .A1(n10), .A2(n629), .ZN(n631) );
  nr02d0 U1115 ( .A1(n10), .A2(n634), .ZN(n636) );
  nr02d0 U1116 ( .A1(n11), .A2(n639), .ZN(n641) );
  nr02d0 U1117 ( .A1(n12), .A2(n644), .ZN(n646) );
  nr02d0 U1118 ( .A1(n11), .A2(n649), .ZN(n651) );
  nr02d0 U1119 ( .A1(n12), .A2(n654), .ZN(n656) );
  nr02d0 U1120 ( .A1(n8), .A2(n659), .ZN(n661) );
  nr02d0 U1121 ( .A1(n9), .A2(n664), .ZN(n666) );
  nr02d0 U1122 ( .A1(n10), .A2(n669), .ZN(n671) );
  inv0d1 U1123 ( .I(s3_op2[17]), .ZN(n674) );
  nr02d0 U1124 ( .A1(n8), .A2(n674), .ZN(n676) );
  inv0d1 U1125 ( .I(s3_op2[18]), .ZN(n679) );
  nr02d0 U1126 ( .A1(n9), .A2(n679), .ZN(n681) );
  inv0d1 U1127 ( .I(s3_op2[19]), .ZN(n684) );
  nr02d0 U1128 ( .A1(n11), .A2(n684), .ZN(n686) );
  inv0d1 U1129 ( .I(s3_op2[20]), .ZN(n689) );
  nr02d0 U1130 ( .A1(n12), .A2(n689), .ZN(n691) );
  inv0d1 U1131 ( .I(s3_op2[21]), .ZN(n694) );
  nr02d0 U1132 ( .A1(n8), .A2(n694), .ZN(n696) );
  inv0d1 U1133 ( .I(s3_op2[22]), .ZN(n699) );
  nr02d0 U1134 ( .A1(n10), .A2(n699), .ZN(n701) );
  inv0d1 U1135 ( .I(s3_op2[23]), .ZN(n704) );
  nr02d0 U1136 ( .A1(n11), .A2(n704), .ZN(n706) );
  inv0d1 U1137 ( .I(s3_op2[24]), .ZN(n709) );
  nr02d0 U1138 ( .A1(n9), .A2(n709), .ZN(n711) );
  inv0d1 U1139 ( .I(s3_op2[25]), .ZN(n714) );
  nr02d0 U1140 ( .A1(n10), .A2(n714), .ZN(n716) );
  inv0d1 U1141 ( .I(s3_op2[26]), .ZN(n719) );
  nr02d0 U1142 ( .A1(n11), .A2(n719), .ZN(n721) );
  nd03d0 U1143 ( .A1(n726), .A2(n725), .A3(n724), .ZN(N893) );
  nd03d0 U1144 ( .A1(n729), .A2(n728), .A3(n727), .ZN(N894) );
  nd03d0 U1145 ( .A1(n732), .A2(n731), .A3(n730), .ZN(N895) );
  nd03d0 U1146 ( .A1(n735), .A2(n734), .A3(n733), .ZN(N896) );
  nd03d0 U1147 ( .A1(n739), .A2(n738), .A3(n737), .ZN(N897) );
  inv0d1 U1148 ( .I(N413), .ZN(n741) );
  inv0d1 U1149 ( .I(n488), .ZN(n851) );
  nd02d1 U1150 ( .A1(N346), .A2(trans3), .ZN(n742) );
  nd03d0 U1151 ( .A1(n744), .A2(n743), .A3(n742), .ZN(N541) );
  inv0d1 U1152 ( .I(N414), .ZN(n745) );
  nr02d0 U1153 ( .A1(n486), .A2(n745), .ZN(n748) );
  inv0d1 U1154 ( .I(s2_op1[1]), .ZN(n746) );
  nr02d0 U1155 ( .A1(n17), .A2(n746), .ZN(n747) );
  nr02d0 U1156 ( .A1(n748), .A2(n747), .ZN(n749) );
  nd02d1 U1157 ( .A1(n750), .A2(n749), .ZN(N542) );
  inv0d1 U1158 ( .I(s2_op1[2]), .ZN(n751) );
  nr02d0 U1159 ( .A1(n468), .A2(n751), .ZN(n753) );
  inv0d1 U1160 ( .I(s2_op1[3]), .ZN(n756) );
  nr02d0 U1161 ( .A1(n470), .A2(n756), .ZN(n758) );
  inv0d1 U1162 ( .I(s2_op1[4]), .ZN(n761) );
  nr02d0 U1163 ( .A1(n471), .A2(n761), .ZN(n763) );
  nd03d0 U1164 ( .A1(n768), .A2(n767), .A3(n766), .ZN(N546) );
  nd03d0 U1165 ( .A1(n771), .A2(n770), .A3(n769), .ZN(N547) );
  nd03d0 U1166 ( .A1(n774), .A2(n773), .A3(n772), .ZN(N548) );
  nd03d0 U1167 ( .A1(n777), .A2(n776), .A3(n775), .ZN(N549) );
  nd03d0 U1168 ( .A1(n780), .A2(n779), .A3(n778), .ZN(N550) );
  nd03d0 U1169 ( .A1(n783), .A2(n782), .A3(n781), .ZN(N551) );
  nd03d0 U1170 ( .A1(n786), .A2(n785), .A3(n784), .ZN(N552) );
  nd03d0 U1171 ( .A1(n789), .A2(n788), .A3(n787), .ZN(N553) );
  nd03d0 U1172 ( .A1(n792), .A2(n791), .A3(n790), .ZN(N554) );
  nd03d0 U1173 ( .A1(n795), .A2(n794), .A3(n793), .ZN(N555) );
  nd03d0 U1174 ( .A1(n798), .A2(n797), .A3(n796), .ZN(N556) );
  nd03d0 U1175 ( .A1(n801), .A2(n800), .A3(n799), .ZN(N557) );
  nd03d0 U1176 ( .A1(n804), .A2(n803), .A3(n802), .ZN(N558) );
  nd03d0 U1177 ( .A1(n807), .A2(n806), .A3(n805), .ZN(N559) );
  nd03d0 U1178 ( .A1(n810), .A2(n809), .A3(n808), .ZN(N560) );
  nd03d0 U1179 ( .A1(n813), .A2(n812), .A3(n811), .ZN(N561) );
  nd03d0 U1180 ( .A1(n816), .A2(n815), .A3(n814), .ZN(N562) );
  nd03d0 U1181 ( .A1(n819), .A2(n818), .A3(n817), .ZN(N563) );
  nd03d0 U1182 ( .A1(n822), .A2(n821), .A3(n820), .ZN(N564) );
  nd03d0 U1183 ( .A1(n825), .A2(n824), .A3(n823), .ZN(N565) );
  nd03d0 U1184 ( .A1(n828), .A2(n827), .A3(n826), .ZN(N566) );
  nd03d0 U1185 ( .A1(n831), .A2(n830), .A3(n829), .ZN(N567) );
  nd03d0 U1186 ( .A1(n834), .A2(n833), .A3(n832), .ZN(N568) );
  nd03d0 U1187 ( .A1(n837), .A2(n836), .A3(n835), .ZN(N569) );
  nd03d0 U1188 ( .A1(n840), .A2(n839), .A3(n838), .ZN(N570) );
  nd03d0 U1189 ( .A1(n843), .A2(n842), .A3(n841), .ZN(N571) );
  nd03d0 U1190 ( .A1(n846), .A2(n845), .A3(n844), .ZN(N572) );
  inv0d1 U1191 ( .I(N445), .ZN(n847) );
  nd02d1 U1192 ( .A1(N378), .A2(trans3), .ZN(n848) );
  nd03d0 U1193 ( .A1(n850), .A2(n849), .A3(n848), .ZN(N573) );
  nd02d1 U1194 ( .A1(N446), .A2(n851), .ZN(n853) );
  nd03d0 U1195 ( .A1(n854), .A2(n853), .A3(n852), .ZN(N574) );
  nd03d0 U1196 ( .A1(n857), .A2(n856), .A3(n855), .ZN(N575) );
  nd03d0 U1197 ( .A1(n860), .A2(n859), .A3(n858), .ZN(N576) );
  nd03d0 U1198 ( .A1(n863), .A2(n862), .A3(n861), .ZN(N577) );
  nd03d0 U1199 ( .A1(n866), .A2(n865), .A3(n864), .ZN(N578) );
  nd03d0 U1200 ( .A1(n869), .A2(n868), .A3(n867), .ZN(N579) );
  nd03d0 U1201 ( .A1(n872), .A2(n871), .A3(n870), .ZN(N580) );
  nd03d0 U1202 ( .A1(n875), .A2(n874), .A3(n873), .ZN(N581) );
  nd03d0 U1203 ( .A1(n878), .A2(n877), .A3(n876), .ZN(N582) );
  nd03d0 U1204 ( .A1(n881), .A2(n880), .A3(n879), .ZN(N583) );
  nd03d0 U1205 ( .A1(n884), .A2(n883), .A3(n882), .ZN(N584) );
  nd03d0 U1206 ( .A1(n887), .A2(n886), .A3(n885), .ZN(N585) );
  nd03d0 U1207 ( .A1(n890), .A2(n889), .A3(n888), .ZN(N586) );
  nd03d0 U1208 ( .A1(n893), .A2(n892), .A3(n891), .ZN(N587) );
  nd03d0 U1209 ( .A1(n896), .A2(n895), .A3(n894), .ZN(N588) );
  nd03d0 U1210 ( .A1(n899), .A2(n898), .A3(n897), .ZN(N589) );
  nd03d0 U1211 ( .A1(n902), .A2(n901), .A3(n900), .ZN(N590) );
  nd03d0 U1212 ( .A1(n905), .A2(n904), .A3(n903), .ZN(N591) );
  nd03d0 U1213 ( .A1(n908), .A2(n907), .A3(n906), .ZN(N592) );
  nd03d0 U1214 ( .A1(n911), .A2(n910), .A3(n909), .ZN(N593) );
  nd03d0 U1215 ( .A1(n914), .A2(n913), .A3(n912), .ZN(N594) );
  nd03d0 U1216 ( .A1(n917), .A2(n916), .A3(n915), .ZN(N595) );
  nd03d0 U1217 ( .A1(n920), .A2(n919), .A3(n918), .ZN(N596) );
  nd03d0 U1218 ( .A1(n923), .A2(n922), .A3(n921), .ZN(N597) );
  nd03d0 U1219 ( .A1(n926), .A2(n925), .A3(n924), .ZN(N598) );
  nd03d0 U1220 ( .A1(n929), .A2(n928), .A3(n927), .ZN(N599) );
  nd03d0 U1221 ( .A1(n932), .A2(n931), .A3(n930), .ZN(N600) );
  nd03d0 U1222 ( .A1(n935), .A2(n934), .A3(n933), .ZN(N601) );
  nd03d0 U1223 ( .A1(n938), .A2(n937), .A3(n936), .ZN(N602) );
  nd03d0 U1224 ( .A1(n941), .A2(n940), .A3(n939), .ZN(N603) );
  nd03d0 U1225 ( .A1(n945), .A2(n944), .A3(n943), .ZN(N604) );
  lanlq1 LOCKUP ( .D(n15), .EN(gclk), .Q(test_so2) );
endmodule


module RISC_CORE ( clk, reset_n, Instrn, Xecutng_Instrn, EndOfInstrn, PSW, 
        Rd_Instr, RESULT_DATA, OUT_VALID, STACK_FULL, test_si1, test_si2, 
        test_se, test_so2 );
  input [31:0] Instrn;
  output [31:0] Xecutng_Instrn;
  output [10:0] PSW;
  output [15:0] RESULT_DATA;
  input clk, reset_n, test_si1, test_si2, test_se;
  output EndOfInstrn, Rd_Instr, OUT_VALID, STACK_FULL, test_so2;
  wire   PushDataIn_11, Latch_Result, Latch_Flags, ALU_Neg, Rd_Oprnd_A,
         Rd_Oprnd_B, Write_RegC, UseData_Imm_Or_RegB, UseData_Imm_Or_ALU,
         Reset_AluRegs, PushEnbl, PopEnbl, n4, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [7:0] Return_Addr;
  wire   [10:8] PopDataOut;
  wire   [15:0] Oprnd_A;
  wire   [15:0] Oprnd_B;
  wire   [15:0] Op_Result;
  wire   [31:0] Crnt_Instrn_2;
  wire   [2:0] Current_State;
  wire   [15:0] RegPort_B;
  wire   [6:0] Addr_A;
  wire   [15:0] RegPort_C;

  ALU I_ALU ( .reset_n(reset_n), .clk(clk), .Oprnd_A(Oprnd_A), .Oprnd_B(
        Oprnd_B), .ALU_OP(Xecutng_Instrn[29:24]), .Latch_Result(Latch_Result), 
        .Latch_Flags(Latch_Flags), .Lachd_Result(Op_Result), .Zro_Flag(
        PushDataIn_11), .Neg_Flag(ALU_Neg), .Carry_Flag(SYNOPSYS_UNCONNECTED_3), .test_se(test_se), .test_si(test_si1) );
  CONTROL I_CONTROL ( .clk(clk), .reset_n(reset_n), .Crnt_Instrn(Crnt_Instrn_2), .Current_State(Current_State), .Neg_Flag(PSW[1]), .Carry_Flag(PSW[0]), 
        .Zro_Flag(PSW[2]), .Latch_Instr(Rd_Instr), .Rd_Oprnd_A(Rd_Oprnd_A), 
        .Rd_Oprnd_B(Rd_Oprnd_B), .Latch_Flags(Latch_Flags), .Latch_Result(
        Latch_Result), .Write_RegC(Write_RegC), .UseData_Imm_Or_RegB(
        UseData_Imm_Or_RegB), .UseData_Imm_Or_ALU(UseData_Imm_Or_ALU), 
        .Reset_AluRegs(Reset_AluRegs), .EndOfInstrn(EndOfInstrn), .PushEnbl(
        PushEnbl), .PopEnbl(PopEnbl), .OUT_VALID(OUT_VALID), .test_se(test_se), 
        .test_si(PushDataIn_11) );
  DATA_PATH I_DATA_PATH ( .clk(clk), .reset_n(reset_n), .Reset_AluRegs(
        Reset_AluRegs), .Rd_Oprnd_A(Rd_Oprnd_A), .Rd_Oprnd_B(Rd_Oprnd_B), 
        .UseData_Imm_Or_RegB(UseData_Imm_Or_RegB), .UseData_Imm_Or_ALU(
        UseData_Imm_Or_ALU), .Latch_Flags(Latch_Flags), .ALU_Zro(PushDataIn_11), .ALU_Neg(ALU_Neg), .ALU_Carry(1'b0), .PSW_Zro(PopDataOut[10]), .PSW_Neg(
        PopDataOut[9]), .PSW_Carry(PopDataOut[8]), .Crnt_Instrn(Crnt_Instrn_2), 
        .RegPort_A(RESULT_DATA), .RegPort_B(RegPort_B), .Op_Result(Op_Result), 
        .Zro_Flag(PSW[2]), .Neg_Flag(PSW[1]), .Carry_Flag(PSW[0]), .Addr_A(
        Addr_A), .Oprnd_A(Oprnd_A), .Oprnd_B(Oprnd_B), .RegPort_C(RegPort_C), 
        .test_se(test_se), .test_si(UseData_Imm_Or_RegB), .test_so(n4) );
  INSTRN_LAT I_INSTRN_LAT ( .clk(clk), .Instrn(Instrn), .Latch_Instr(Rd_Instr), 
        .Crnt_Instrn_1(Xecutng_Instrn), .Crnt_Instrn_2(Crnt_Instrn_2), 
        .test_se(test_se), .test_si1(n4), .test_si2(test_si2) );
  PRGRM_CNT_TOP I_PRGRM_CNT_TOP ( .clk(clk), .reset_n(reset_n), .Crnt_Instrn(
        Crnt_Instrn_2), .Zro_Flag(PSW[2]), .Carry_Flag(PSW[0]), .Neg_Flag(
        PSW[1]), .Return_Addr(Return_Addr), .Current_State(Current_State), 
        .PC(PSW[10:3]), .test_si(Crnt_Instrn_2[31]), .test_se(test_se) );
  REG_FILE I_REG_FILE ( .reset_n(reset_n), .clk(clk), .Addr_A(Addr_A), 
        .Addr_B(Xecutng_Instrn[6:0]), .Addr_C(Xecutng_Instrn[22:16]), 
        .RegPort_C(RegPort_C), .Write_RegC(Write_RegC), .RegPort_A(RESULT_DATA), .RegPort_B(RegPort_B) );
  STACK_TOP I_STACK_TOP ( .reset_n(reset_n), .clk(clk), .PushEnbl(PushEnbl), 
        .PopEnbl(PopEnbl), .PushDataIn({PushDataIn_11, PSW[2:0], PSW[10:3]}), 
        .PopDataOut({SYNOPSYS_UNCONNECTED_4, PopDataOut, Return_Addr}), 
        .STACK_FULL(STACK_FULL), .test_si(Current_State[2]), .test_se(test_se), 
        .test_so(test_so2) );
endmodule


module CONTEXT_MEM ( sys_clk, sys_rst_n, context_en, cmd, pci_data_in, 
        pci_context_data );
  input [7:0] cmd;
  input [31:0] pci_data_in;
  output [31:0] pci_context_data;
  input sys_clk, sys_rst_n, context_en;


  bufbd1 U1 ( .I(pci_data_in[31]), .Z(pci_context_data[31]) );
  bufbd1 U2 ( .I(pci_data_in[30]), .Z(pci_context_data[30]) );
  bufbd1 U3 ( .I(pci_data_in[29]), .Z(pci_context_data[29]) );
  bufbd1 U4 ( .I(pci_data_in[28]), .Z(pci_context_data[28]) );
  bufbd1 U5 ( .I(pci_data_in[27]), .Z(pci_context_data[27]) );
  bufbd1 U6 ( .I(pci_data_in[26]), .Z(pci_context_data[26]) );
  bufbd1 U7 ( .I(pci_data_in[25]), .Z(pci_context_data[25]) );
  bufbd1 U8 ( .I(pci_data_in[24]), .Z(pci_context_data[24]) );
  bufbd1 U9 ( .I(pci_data_in[23]), .Z(pci_context_data[23]) );
  bufbd1 U10 ( .I(pci_data_in[22]), .Z(pci_context_data[22]) );
  bufbd1 U11 ( .I(pci_data_in[21]), .Z(pci_context_data[21]) );
  bufbd1 U12 ( .I(pci_data_in[20]), .Z(pci_context_data[20]) );
  bufbd1 U13 ( .I(pci_data_in[19]), .Z(pci_context_data[19]) );
  bufbd1 U14 ( .I(pci_data_in[18]), .Z(pci_context_data[18]) );
  bufbd1 U15 ( .I(pci_data_in[17]), .Z(pci_context_data[17]) );
  bufbd1 U16 ( .I(pci_data_in[16]), .Z(pci_context_data[16]) );
  bufbd1 U17 ( .I(pci_data_in[15]), .Z(pci_context_data[15]) );
  bufbd1 U18 ( .I(pci_data_in[14]), .Z(pci_context_data[14]) );
  bufbd1 U19 ( .I(pci_data_in[13]), .Z(pci_context_data[13]) );
  bufbd1 U20 ( .I(pci_data_in[12]), .Z(pci_context_data[12]) );
  bufbd1 U21 ( .I(pci_data_in[11]), .Z(pci_context_data[11]) );
  bufbd1 U22 ( .I(pci_data_in[10]), .Z(pci_context_data[10]) );
  bufbd1 U23 ( .I(pci_data_in[9]), .Z(pci_context_data[9]) );
  bufbd1 U24 ( .I(pci_data_in[8]), .Z(pci_context_data[8]) );
  bufbd1 U25 ( .I(pci_data_in[7]), .Z(pci_context_data[7]) );
  bufbd1 U26 ( .I(pci_data_in[6]), .Z(pci_context_data[6]) );
  bufbd1 U27 ( .I(pci_data_in[5]), .Z(pci_context_data[5]) );
  bufbd1 U28 ( .I(pci_data_in[4]), .Z(pci_context_data[4]) );
  bufbd1 U29 ( .I(pci_data_in[3]), .Z(pci_context_data[3]) );
  bufbd1 U30 ( .I(pci_data_in[2]), .Z(pci_context_data[2]) );
  bufbd1 U31 ( .I(pci_data_in[1]), .Z(pci_context_data[1]) );
  bufbd1 U32 ( .I(pci_data_in[0]), .Z(pci_context_data[0]) );
endmodule


module PARSER ( sys_clk, pclk, sys_rst_n, pcmd, pcmd_valid, pcmd_out, 
        pcmd_out_valid, blender_op, blender_clk_en, context_en, context_cmd, 
        fifo_read_pop, fifo_read_empty, fifo_write_push, fifo_write_full, 
        risc_Instrn_lo, risc_Xecutng_Instrn_lo, pci_w_mux_select, 
        sd_w_mux_select, parser_sd_rfifo_pop, sd_rfifo_parser_empty, 
        parser_sd_wfifo_push, sd_wfifo_parser_full, test_se, test_si1, 
        test_si2, test_so2, test_so1 );
  input [3:0] pcmd;
  output [3:0] pcmd_out;
  output [3:0] blender_op;
  output [7:0] context_cmd;
  output [7:0] risc_Instrn_lo;
  input [15:0] risc_Xecutng_Instrn_lo;
  output [1:0] pci_w_mux_select;
  output [1:0] sd_w_mux_select;
  input sys_clk, pclk, sys_rst_n, pcmd_valid, fifo_read_empty, fifo_write_full,
         sd_rfifo_parser_empty, sd_wfifo_parser_full, test_se, test_si1,
         test_si2;
  output pcmd_out_valid, blender_clk_en, context_en, fifo_read_pop,
         fifo_write_push, parser_sd_rfifo_pop, parser_sd_wfifo_push, test_so2,
         test_so1;
  wire   r_pcmd_valid, i_pcmd_out_valid, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N31, N32, N33, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N111, N112, N113, N114,
         n48, n50, n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74,
         n76, n78, n81, n84, n87, n90, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n1, n2, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175;
  wire   [3:0] r_pcmd;
  wire   [3:0] sync_pcmd;
  wire   [3:0] sync_pcmd_out;
  wire   [3:0] i_pcmd_out;
  wire   [19:0] i_reg;

  sdnrn1 r_pcmd_reg_2_ ( .D(sync_pcmd[2]), .SD(n87), .SC(test_se), .CP(sys_clk), .QN(n90) );
  sdnrn1 r_pcmd_reg_1_ ( .D(sync_pcmd[1]), .SD(n84), .SC(test_se), .CP(sys_clk), .QN(n87) );
  sdnrn1 r_pcmd_reg_0_ ( .D(sync_pcmd[0]), .SD(pci_w_mux_select[1]), .SC(
        test_se), .CP(sys_clk), .QN(n84) );
  sdnrn1 r_pcmd_valid_reg ( .D(test_so1), .SD(r_pcmd[3]), .SC(test_se), .CP(
        sys_clk), .QN(n81) );
  sdnrn1 i_reg_reg_19_ ( .D(N28), .SD(n105), .SC(test_se), .CP(sys_clk), .QN(
        n78) );
  sdnrn1 i_reg_reg_18_ ( .D(N27), .SD(n108), .SC(test_se), .CP(sys_clk), .QN(
        n76) );
  sdnrn1 i_reg_reg_17_ ( .D(N26), .SD(n111), .SC(test_se), .CP(sys_clk), .QN(
        n74) );
  sdnrn1 i_reg_reg_16_ ( .D(N25), .SD(n114), .SC(test_se), .CP(sys_clk), .QN(
        n72) );
  sdnrn1 i_reg_reg_15_ ( .D(N24), .SD(n117), .SC(test_se), .CP(sys_clk), .QN(
        n70) );
  sdnrn1 i_reg_reg_14_ ( .D(N23), .SD(n120), .SC(test_se), .CP(sys_clk), .QN(
        n68) );
  sdnrn1 i_reg_reg_13_ ( .D(N22), .SD(n123), .SC(test_se), .CP(sys_clk), .QN(
        n66) );
  sdnrn1 i_reg_reg_12_ ( .D(N21), .SD(n127), .SC(test_se), .CP(sys_clk), .QN(
        n64) );
  sdnrn1 i_reg_reg_11_ ( .D(N20), .SD(n128), .SC(test_se), .CP(sys_clk), .QN(
        n62) );
  sdnrn1 i_reg_reg_10_ ( .D(N19), .SD(n132), .SC(test_se), .CP(sys_clk), .QN(
        n60) );
  sdnrn1 i_reg_reg_9_ ( .D(N18), .SD(n136), .SC(test_se), .CP(sys_clk), .QN(
        n58) );
  sdnrn1 i_reg_reg_8_ ( .D(N17), .SD(n138), .SC(test_se), .CP(sys_clk), .QN(
        n56) );
  sdnrn1 i_reg_reg_7_ ( .D(N16), .SD(n140), .SC(test_se), .CP(sys_clk), .QN(
        n54) );
  sdnrn1 i_reg_reg_6_ ( .D(N15), .SD(n142), .SC(test_se), .CP(sys_clk), .QN(
        n52) );
  sdnrn1 i_reg_reg_5_ ( .D(N14), .SD(n144), .SC(test_se), .CP(sys_clk), .QN(
        n50) );
  sdnrn1 i_reg_reg_4_ ( .D(N13), .SD(i_reg[3]), .SC(test_se), .CP(sys_clk), 
        .QN(n48) );
  an02d1 U94 ( .A1(risc_Instrn_lo[0]), .A2(context_cmd[0]), .Z(context_en) );
  an02d1 U113 ( .A1(n147), .A2(r_pcmd_valid), .Z(n135) );
  an04d1 U120 ( .A1(r_pcmd[3]), .A2(r_pcmd[1]), .A3(n161), .A4(n150), .Z(n149)
         );
  aor21d1 U126 ( .B1(i_reg[18]), .B2(n81), .A(n169), .Z(N99) );
  aor21d1 U127 ( .B1(i_reg[17]), .B2(n81), .A(n169), .Z(N98) );
  aor21d1 U128 ( .B1(i_reg[16]), .B2(n81), .A(n167), .Z(N97) );
  aor211d1 U129 ( .C1(i_reg[15]), .C2(n81), .A(n96), .B(n97), .Z(N96) );
  aor222d1 U130 ( .A1(i_reg[19]), .A2(n98), .B1(n99), .B2(i_reg[17]), .C1(n100), .C2(i_reg[16]), .Z(n97) );
  aor22d1 U131 ( .A1(n169), .A2(n101), .B1(n102), .B2(i_reg[18]), .Z(n96) );
  aor211d1 U132 ( .C1(i_reg[14]), .C2(n81), .A(n103), .B(n104), .Z(N95) );
  aor222d1 U133 ( .A1(n98), .A2(i_reg[18]), .B1(n99), .B2(i_reg[16]), .C1(
        i_reg[15]), .C2(n100), .Z(n104) );
  aor22d1 U134 ( .A1(n169), .A2(n105), .B1(n102), .B2(i_reg[17]), .Z(n103) );
  aor211d1 U135 ( .C1(i_reg[13]), .C2(n81), .A(n106), .B(n107), .Z(N94) );
  aor222d1 U136 ( .A1(n98), .A2(i_reg[17]), .B1(i_reg[15]), .B2(n99), .C1(
        i_reg[14]), .C2(n100), .Z(n107) );
  aor22d1 U137 ( .A1(n167), .A2(n108), .B1(n102), .B2(i_reg[16]), .Z(n106) );
  aor211d1 U138 ( .C1(i_reg[12]), .C2(n81), .A(n109), .B(n110), .Z(N93) );
  aor222d1 U139 ( .A1(n98), .A2(i_reg[16]), .B1(i_reg[14]), .B2(n99), .C1(
        i_reg[13]), .C2(n100), .Z(n110) );
  aor22d1 U140 ( .A1(n167), .A2(n111), .B1(i_reg[15]), .B2(n102), .Z(n109) );
  aor211d1 U141 ( .C1(i_reg[11]), .C2(n81), .A(n112), .B(n113), .Z(N92) );
  aor222d1 U142 ( .A1(i_reg[15]), .A2(n98), .B1(i_reg[13]), .B2(n99), .C1(
        i_reg[12]), .C2(n100), .Z(n113) );
  aor22d1 U143 ( .A1(n169), .A2(n114), .B1(i_reg[14]), .B2(n102), .Z(n112) );
  aor211d1 U144 ( .C1(i_reg[10]), .C2(n81), .A(n115), .B(n116), .Z(N91) );
  aor222d1 U145 ( .A1(i_reg[14]), .A2(n98), .B1(i_reg[12]), .B2(n99), .C1(
        i_reg[11]), .C2(n100), .Z(n116) );
  aor22d1 U146 ( .A1(n169), .A2(n117), .B1(i_reg[13]), .B2(n102), .Z(n115) );
  aor211d1 U147 ( .C1(i_reg[9]), .C2(n81), .A(n118), .B(n119), .Z(N90) );
  aor222d1 U148 ( .A1(i_reg[13]), .A2(n98), .B1(i_reg[11]), .B2(n99), .C1(
        i_reg[10]), .C2(n100), .Z(n119) );
  aor22d1 U149 ( .A1(n167), .A2(n120), .B1(i_reg[12]), .B2(n102), .Z(n118) );
  xr02d1 U150 ( .A1(sd_wfifo_parser_full), .A2(sd_rfifo_parser_empty), .Z(N9)
         );
  aor211d1 U151 ( .C1(i_reg[8]), .C2(n81), .A(n121), .B(n122), .Z(N89) );
  aor222d1 U152 ( .A1(i_reg[12]), .A2(n98), .B1(i_reg[10]), .B2(n99), .C1(
        i_reg[9]), .C2(n100), .Z(n122) );
  aor22d1 U153 ( .A1(n167), .A2(n123), .B1(i_reg[11]), .B2(n102), .Z(n121) );
  aor211d1 U154 ( .C1(i_reg[7]), .C2(n81), .A(n124), .B(n125), .Z(N88) );
  aor222d1 U155 ( .A1(i_reg[11]), .A2(n98), .B1(i_reg[9]), .B2(n99), .C1(
        i_reg[8]), .C2(n100), .Z(n125) );
  aor22d1 U157 ( .A1(n169), .A2(n127), .B1(i_reg[10]), .B2(n102), .Z(n124) );
  aor221d1 U158 ( .B1(i_reg[9]), .B2(n102), .C1(n169), .C2(n128), .A(n129), 
        .Z(N87) );
  aor222d1 U159 ( .A1(i_reg[10]), .A2(n98), .B1(i_reg[6]), .B2(n130), .C1(
        i_reg[7]), .C2(n100), .Z(n129) );
  aor221d1 U160 ( .B1(i_reg[8]), .B2(n102), .C1(n167), .C2(n132), .A(n133), 
        .Z(N86) );
  aor222d1 U161 ( .A1(i_reg[5]), .A2(n134), .B1(n135), .B2(i_reg[9]), .C1(
        i_reg[6]), .C2(n100), .Z(n133) );
  aor221d1 U162 ( .B1(i_reg[7]), .B2(n102), .C1(n167), .C2(n136), .A(n137), 
        .Z(N85) );
  aor222d1 U163 ( .A1(i_reg[4]), .A2(n134), .B1(n135), .B2(i_reg[8]), .C1(
        i_reg[5]), .C2(n100), .Z(n137) );
  aor221d1 U164 ( .B1(i_reg[6]), .B2(n102), .C1(n169), .C2(n138), .A(n139), 
        .Z(N84) );
  aor222d1 U165 ( .A1(i_reg[3]), .A2(n134), .B1(n135), .B2(i_reg[7]), .C1(
        i_reg[4]), .C2(n100), .Z(n139) );
  aor221d1 U166 ( .B1(i_reg[5]), .B2(n102), .C1(n169), .C2(n140), .A(n141), 
        .Z(N83) );
  aor222d1 U167 ( .A1(i_reg[2]), .A2(n134), .B1(n135), .B2(i_reg[6]), .C1(
        i_reg[3]), .C2(n100), .Z(n141) );
  aor221d1 U168 ( .B1(i_reg[4]), .B2(n102), .C1(n167), .C2(n142), .A(n143), 
        .Z(N82) );
  aor222d1 U169 ( .A1(i_reg[1]), .A2(n134), .B1(i_reg[5]), .B2(n135), .C1(
        i_reg[2]), .C2(n100), .Z(n143) );
  aor221d1 U170 ( .B1(i_reg[3]), .B2(n102), .C1(n167), .C2(n144), .A(n145), 
        .Z(N81) );
  aor222d1 U171 ( .A1(i_reg[0]), .A2(n134), .B1(i_reg[4]), .B2(n135), .C1(
        i_reg[1]), .C2(n100), .Z(n145) );
  nd03d0 U172 ( .A1(n148), .A2(n126), .A3(r_pcmd_valid), .ZN(n134) );
  nr02d0 U173 ( .A1(n150), .A2(n81), .ZN(N8) );
  xr02d1 U174 ( .A1(i_reg[17]), .A2(i_reg[13]), .Z(N33) );
  xr02d1 U175 ( .A1(sd_wfifo_parser_full), .A2(fifo_read_empty), .Z(N28) );
  xr02d1 U176 ( .A1(fifo_write_full), .A2(fifo_read_empty), .Z(N27) );
  xr02d1 U177 ( .A1(risc_Xecutng_Instrn_lo[15]), .A2(fifo_write_full), .Z(N26)
         );
  xr02d1 U178 ( .A1(risc_Xecutng_Instrn_lo[15]), .A2(
        risc_Xecutng_Instrn_lo[14]), .Z(N25) );
  xr02d1 U179 ( .A1(risc_Xecutng_Instrn_lo[14]), .A2(
        risc_Xecutng_Instrn_lo[13]), .Z(N24) );
  xr02d1 U180 ( .A1(risc_Xecutng_Instrn_lo[13]), .A2(
        risc_Xecutng_Instrn_lo[12]), .Z(N23) );
  xr02d1 U181 ( .A1(risc_Xecutng_Instrn_lo[12]), .A2(
        risc_Xecutng_Instrn_lo[11]), .Z(N22) );
  xr02d1 U182 ( .A1(risc_Xecutng_Instrn_lo[11]), .A2(
        risc_Xecutng_Instrn_lo[10]), .Z(N21) );
  xr02d1 U183 ( .A1(risc_Xecutng_Instrn_lo[9]), .A2(risc_Xecutng_Instrn_lo[10]), .Z(N20) );
  xr02d1 U184 ( .A1(risc_Xecutng_Instrn_lo[9]), .A2(risc_Xecutng_Instrn_lo[8]), 
        .Z(N19) );
  xr02d1 U185 ( .A1(risc_Xecutng_Instrn_lo[8]), .A2(risc_Xecutng_Instrn_lo[7]), 
        .Z(N18) );
  xr02d1 U186 ( .A1(risc_Xecutng_Instrn_lo[7]), .A2(risc_Xecutng_Instrn_lo[6]), 
        .Z(N17) );
  xr02d1 U187 ( .A1(risc_Xecutng_Instrn_lo[6]), .A2(risc_Xecutng_Instrn_lo[5]), 
        .Z(N16) );
  xr02d1 U188 ( .A1(risc_Xecutng_Instrn_lo[5]), .A2(risc_Xecutng_Instrn_lo[4]), 
        .Z(N15) );
  xr02d1 U189 ( .A1(risc_Xecutng_Instrn_lo[4]), .A2(risc_Xecutng_Instrn_lo[3]), 
        .Z(N14) );
  xr02d1 U190 ( .A1(risc_Xecutng_Instrn_lo[3]), .A2(risc_Xecutng_Instrn_lo[2]), 
        .Z(N13) );
  xr02d1 U191 ( .A1(risc_Xecutng_Instrn_lo[2]), .A2(risc_Xecutng_Instrn_lo[1]), 
        .Z(N12) );
  nd23d1 U192 ( .A1(n151), .A2(n152), .A3(n153), .ZN(N114) );
  nr02d0 U193 ( .A1(n151), .A2(n154), .ZN(N113) );
  nr04d0 U194 ( .A1(n155), .A2(n156), .A3(risc_Xecutng_Instrn_lo[1]), .A4(
        sd_rfifo_parser_empty), .ZN(n151) );
  nd23d1 U195 ( .A1(n154), .A2(n157), .A3(n153), .ZN(N112) );
  nd04d0 U196 ( .A1(risc_Xecutng_Instrn_lo[0]), .A2(risc_Xecutng_Instrn_lo[1]), 
        .A3(sd_rfifo_parser_empty), .A4(sd_wfifo_parser_full), .ZN(n153) );
  nr04d0 U197 ( .A1(n158), .A2(n156), .A3(risc_Xecutng_Instrn_lo[0]), .A4(
        sd_rfifo_parser_empty), .ZN(n154) );
  nr02d0 U198 ( .A1(n152), .A2(n157), .ZN(N111) );
  nr04d0 U199 ( .A1(n158), .A2(n159), .A3(risc_Xecutng_Instrn_lo[0]), .A4(
        sd_wfifo_parser_full), .ZN(n157) );
  nr04d0 U200 ( .A1(n155), .A2(n159), .A3(risc_Xecutng_Instrn_lo[1]), .A4(
        sd_wfifo_parser_full), .ZN(n152) );
  xr02d1 U201 ( .A1(risc_Xecutng_Instrn_lo[1]), .A2(risc_Xecutng_Instrn_lo[0]), 
        .Z(N11) );
  aor21d1 U202 ( .B1(i_reg[19]), .B2(n81), .A(n167), .Z(N100) );
  nr03d0 U203 ( .A1(n81), .A2(n131), .A3(n160), .ZN(n95) );
  nd23d1 U204 ( .A1(n146), .A2(n149), .A3(n126), .ZN(n160) );
  nd04d0 U205 ( .A1(r_pcmd[2]), .A2(r_pcmd[3]), .A3(n161), .A4(n162), .ZN(n126) );
  nr04d0 U206 ( .A1(n161), .A2(n162), .A3(r_pcmd[2]), .A4(r_pcmd[3]), .ZN(n146) );
  nd04d0 U207 ( .A1(r_pcmd[0]), .A2(r_pcmd[3]), .A3(n162), .A4(n150), .ZN(n148) );
  nr04d0 U208 ( .A1(n161), .A2(n150), .A3(r_pcmd[1]), .A4(r_pcmd[3]), .ZN(n147) );
  xr02d1 U209 ( .A1(sd_rfifo_parser_empty), .A2(risc_Xecutng_Instrn_lo[0]), 
        .Z(N10) );
  sdcrq1 out_bus_reg_8_ ( .D(N89), .SD(risc_Instrn_lo[7]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(blender_op[0]) );
  sdcrq1 out_bus_reg_9_ ( .D(N90), .SD(context_cmd[0]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(blender_op[1]) );
  sdcrq1 out_bus_reg_10_ ( .D(N91), .SD(context_cmd[1]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(blender_op[2]) );
  sdcrq1 out_bus_reg_11_ ( .D(N92), .SD(context_cmd[2]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(blender_op[3]) );
  sdnrq1 r_pcmd_out_valid_reg ( .D(test_so2), .SD(pcmd_out[3]), .SC(test_se), 
        .CP(pclk), .Q(pcmd_out_valid) );
  sdnrq1 r_pcmd_out_reg_0_ ( .D(sync_pcmd_out[0]), .SD(test_si2), .SC(test_se), 
        .CP(pclk), .Q(pcmd_out[0]) );
  sdnrq1 r_pcmd_out_reg_2_ ( .D(sync_pcmd_out[2]), .SD(pcmd_out[1]), .SC(
        test_se), .CP(pclk), .Q(pcmd_out[2]) );
  sdnrq1 r_pcmd_out_reg_1_ ( .D(sync_pcmd_out[1]), .SD(pcmd_out[0]), .SC(
        test_se), .CP(pclk), .Q(pcmd_out[1]) );
  sdnrq1 r_pcmd_out_reg_3_ ( .D(sync_pcmd_out[3]), .SD(pcmd_out[2]), .SC(
        test_se), .CP(pclk), .Q(pcmd_out[3]) );
  sdcrq1 pci_w_mux_select_reg_1_ ( .D(N112), .SD(pci_w_mux_select[0]), .SC(
        test_se), .CP(sys_clk), .CDN(sys_rst_n), .Q(pci_w_mux_select[1]) );
  sdnrq1 i_reg_reg_3_ ( .D(N12), .SD(i_reg[2]), .SC(test_se), .CP(sys_clk), 
        .Q(i_reg[3]) );
  sdcrq1 pci_w_mux_select_reg_0_ ( .D(N111), .SD(context_cmd[7]), .SC(test_se), 
        .CP(sys_clk), .CDN(sys_rst_n), .Q(pci_w_mux_select[0]) );
  sdnrq1 i_reg_reg_2_ ( .D(N11), .SD(i_reg[1]), .SC(test_se), .CP(sys_clk), 
        .Q(i_reg[2]) );
  sdnrq1 r_pcmd_reg_3_ ( .D(sync_pcmd[3]), .SD(n90), .SC(test_se), .CP(sys_clk), .Q(r_pcmd[3]) );
  sdnrq1 i_reg_reg_1_ ( .D(N10), .SD(i_reg[0]), .SC(test_se), .CP(sys_clk), 
        .Q(i_reg[1]) );
  sdnrq1 i_reg_reg_0_ ( .D(N9), .SD(i_pcmd_out_valid), .SC(test_se), .CP(
        sys_clk), .Q(i_reg[0]) );
  sdcrq1 sd_w_mux_select_reg_1_ ( .D(N114), .SD(sd_w_mux_select[0]), .SC(
        test_se), .CP(sys_clk), .CDN(sys_rst_n), .Q(sd_w_mux_select[1]) );
  sdcrq1 sd_w_mux_select_reg_0_ ( .D(N113), .SD(n81), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(sd_w_mux_select[0]) );
  sdcrq1 out_bus_reg_15_ ( .D(N96), .SD(parser_sd_rfifo_pop), .SC(test_se), 
        .CP(sys_clk), .CDN(sys_rst_n), .Q(parser_sd_wfifo_push) );
  sdcrq1 out_bus_reg_14_ ( .D(N95), .SD(fifo_write_push), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(parser_sd_rfifo_pop) );
  sdcrq1 out_bus_reg_12_ ( .D(N93), .SD(context_cmd[3]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(fifo_read_pop) );
  sdcrq1 out_bus_reg_13_ ( .D(N94), .SD(fifo_read_pop), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(fifo_write_push) );
  sdcrq1 i_pcmd_out_reg_3_ ( .D(N32), .SD(i_pcmd_out[2]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(i_pcmd_out[3]) );
  sdcrq1 i_pcmd_out_reg_2_ ( .D(N31), .SD(i_pcmd_out[1]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(i_pcmd_out[2]) );
  sdcrq1 i_pcmd_out_reg_1_ ( .D(n1), .SD(i_pcmd_out[0]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(i_pcmd_out[1]) );
  sdcrq1 i_pcmd_out_reg_0_ ( .D(N29), .SD(blender_clk_en), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(i_pcmd_out[0]) );
  sdcrq1 out_bus_reg_3_ ( .D(N84), .SD(risc_Instrn_lo[2]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[3]) );
  sdcrq1 out_bus_reg_2_ ( .D(N83), .SD(risc_Instrn_lo[1]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[2]) );
  sdcrq1 out_bus_reg_1_ ( .D(N82), .SD(risc_Instrn_lo[0]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[1]) );
  sdcrq1 out_bus_reg_0_ ( .D(N81), .SD(n101), .SC(test_se), .CP(sys_clk), 
        .CDN(sys_rst_n), .Q(risc_Instrn_lo[0]) );
  sdcrq1 out_bus_reg_19_ ( .D(N100), .SD(context_cmd[6]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(context_cmd[7]) );
  sdcrq1 out_bus_reg_18_ ( .D(N99), .SD(context_cmd[5]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(context_cmd[6]) );
  sdcrq1 out_bus_reg_17_ ( .D(N98), .SD(context_cmd[4]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(context_cmd[5]) );
  sdcrq1 out_bus_reg_16_ ( .D(N97), .SD(parser_sd_wfifo_push), .SC(test_se), 
        .CP(sys_clk), .CDN(sys_rst_n), .Q(context_cmd[4]) );
  sdcrq1 i_pcmd_out_valid_reg ( .D(N33), .SD(i_pcmd_out[3]), .SC(test_se), 
        .CP(sys_clk), .CDN(sys_rst_n), .Q(i_pcmd_out_valid) );
  sdcrq1 out_bus_reg_7_ ( .D(N88), .SD(risc_Instrn_lo[6]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[7]) );
  sdcrq1 out_bus_reg_6_ ( .D(N87), .SD(risc_Instrn_lo[5]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[6]) );
  sdcrq1 out_bus_reg_5_ ( .D(N86), .SD(risc_Instrn_lo[4]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[5]) );
  sdcrq1 out_bus_reg_4_ ( .D(N85), .SD(risc_Instrn_lo[3]), .SC(test_se), .CP(
        sys_clk), .CDN(sys_rst_n), .Q(risc_Instrn_lo[4]) );
  sdcrq1 blender_clk_en_reg ( .D(N8), .SD(test_si1), .SC(test_se), .CP(sys_clk), .CDN(sys_rst_n), .Q(blender_clk_en) );
  sdnrq1 sync_pcmd_out_valid_reg ( .D(i_pcmd_out_valid), .SD(sync_pcmd_out[3]), 
        .SC(test_se), .CP(pclk), .Q(test_so2) );
  sdnrq1 sync_pcmd_out_reg_3_ ( .D(i_pcmd_out[3]), .SD(sync_pcmd_out[2]), .SC(
        test_se), .CP(pclk), .Q(sync_pcmd_out[3]) );
  sdnrq1 sync_pcmd_out_reg_2_ ( .D(i_pcmd_out[2]), .SD(sync_pcmd_out[1]), .SC(
        test_se), .CP(pclk), .Q(sync_pcmd_out[2]) );
  sdnrq1 sync_pcmd_out_reg_1_ ( .D(i_pcmd_out[1]), .SD(sync_pcmd_out[0]), .SC(
        test_se), .CP(pclk), .Q(sync_pcmd_out[1]) );
  sdnrq1 sync_pcmd_out_reg_0_ ( .D(i_pcmd_out[0]), .SD(pcmd_out_valid), .SC(
        test_se), .CP(pclk), .Q(sync_pcmd_out[0]) );
  sdnrq1 sync_pcmd_reg_3_ ( .D(pcmd[3]), .SD(sync_pcmd[2]), .SC(test_se), .CP(
        sys_clk), .Q(sync_pcmd[3]) );
  sdnrq1 sync_pcmd_reg_2_ ( .D(pcmd[2]), .SD(sync_pcmd[1]), .SC(test_se), .CP(
        sys_clk), .Q(sync_pcmd[2]) );
  sdnrq1 sync_pcmd_reg_1_ ( .D(pcmd[1]), .SD(sync_pcmd[0]), .SC(test_se), .CP(
        sys_clk), .Q(sync_pcmd[1]) );
  sdnrq1 sync_pcmd_reg_0_ ( .D(pcmd[0]), .SD(sd_w_mux_select[1]), .SC(test_se), 
        .CP(sys_clk), .Q(sync_pcmd[0]) );
  sdnrq1 sync_pcmd_valid_reg ( .D(pcmd_valid), .SD(sync_pcmd[3]), .SC(test_se), 
        .CP(sys_clk), .Q(test_so1) );
  bufbd1 U4 ( .I(blender_op[0]), .Z(context_cmd[0]) );
  bufbd1 U48 ( .I(blender_op[2]), .Z(context_cmd[2]) );
  bufbd1 U50 ( .I(blender_op[1]), .Z(context_cmd[1]) );
  bufbd1 U52 ( .I(blender_op[3]), .Z(context_cmd[3]) );
  inv0d1 U54 ( .I(n168), .ZN(n169) );
  inv0d1 U56 ( .I(n95), .ZN(n168) );
  inv0d1 U58 ( .I(n166), .ZN(n167) );
  inv0d1 U60 ( .I(n165), .ZN(n166) );
  inv0d1 U62 ( .I(sd_rfifo_parser_empty), .ZN(n159) );
  inv0d1 U64 ( .I(i_reg[15]), .ZN(n114) );
  inv0d1 U66 ( .I(i_reg[14]), .ZN(n117) );
  inv0d1 U68 ( .I(i_reg[11]), .ZN(n127) );
  inv0d1 U70 ( .I(i_reg[18]), .ZN(n105) );
  inv0d1 U72 ( .I(i_reg[19]), .ZN(n101) );
  inv0d1 U74 ( .I(i_reg[8]), .ZN(n136) );
  inv0d1 U76 ( .I(i_reg[9]), .ZN(n132) );
  inv0d1 U78 ( .I(i_reg[13]), .ZN(n120) );
  inv0d1 U81 ( .I(i_reg[12]), .ZN(n123) );
  inv0d1 U84 ( .I(i_reg[16]), .ZN(n111) );
  inv0d1 U87 ( .I(i_reg[17]), .ZN(n108) );
  inv0d1 U90 ( .I(r_pcmd[0]), .ZN(n161) );
  inv0d1 U95 ( .I(r_pcmd[1]), .ZN(n162) );
  an02d1 U96 ( .A1(n146), .A2(r_pcmd_valid), .Z(n100) );
  an02d1 U97 ( .A1(n149), .A2(r_pcmd_valid), .Z(n102) );
  nd12d0 U98 ( .A1(n147), .A2(n148), .ZN(n131) );
  an02d1 U99 ( .A1(r_pcmd_valid), .A2(n131), .Z(n98) );
  nr02d0 U100 ( .A1(n126), .A2(n81), .ZN(n99) );
  inv0d1 U101 ( .I(i_reg[10]), .ZN(n128) );
  nd02d1 U102 ( .A1(r_pcmd_valid), .A2(n126), .ZN(n130) );
  inv0d1 U103 ( .I(i_reg[9]), .ZN(n171) );
  inv0d1 U104 ( .I(r_pcmd[2]), .ZN(n150) );
  inv0d1 U105 ( .I(n174), .ZN(n172) );
  inv0d1 U106 ( .I(risc_Xecutng_Instrn_lo[1]), .ZN(n158) );
  inv0d1 U107 ( .I(risc_Xecutng_Instrn_lo[0]), .ZN(n155) );
  inv0d1 U108 ( .I(i_reg[4]), .ZN(n144) );
  inv0d1 U109 ( .I(i_reg[5]), .ZN(n142) );
  inv0d1 U110 ( .I(i_reg[6]), .ZN(n140) );
  inv0d1 U111 ( .I(i_reg[7]), .ZN(n138) );
  inv0d1 U112 ( .I(n87), .ZN(r_pcmd[1]) );
  inv0d1 U114 ( .I(n90), .ZN(r_pcmd[2]) );
  inv0d1 U115 ( .I(n84), .ZN(r_pcmd[0]) );
  inv0d1 U116 ( .I(n81), .ZN(r_pcmd_valid) );
  inv0d1 U117 ( .I(n54), .ZN(i_reg[7]) );
  inv0d1 U118 ( .I(n58), .ZN(i_reg[9]) );
  inv0d1 U119 ( .I(n60), .ZN(i_reg[10]) );
  inv0d1 U121 ( .I(n56), .ZN(i_reg[8]) );
  inv0d1 U122 ( .I(n66), .ZN(i_reg[13]) );
  inv0d1 U123 ( .I(n74), .ZN(i_reg[17]) );
  inv0d1 U124 ( .I(n72), .ZN(i_reg[16]) );
  inv0d1 U125 ( .I(n68), .ZN(i_reg[14]) );
  inv0d1 U156 ( .I(n64), .ZN(i_reg[12]) );
  inv0d1 U210 ( .I(n62), .ZN(i_reg[11]) );
  inv0d1 U211 ( .I(n70), .ZN(i_reg[15]) );
  inv0d1 U212 ( .I(sd_wfifo_parser_full), .ZN(n156) );
  inv0d1 U213 ( .I(n52), .ZN(i_reg[6]) );
  inv0d1 U214 ( .I(n48), .ZN(i_reg[4]) );
  inv0d1 U215 ( .I(n50), .ZN(i_reg[5]) );
  inv0d1 U216 ( .I(n76), .ZN(i_reg[18]) );
  inv0d1 U217 ( .I(n78), .ZN(i_reg[19]) );
  xr03d1 U218 ( .A1(i_reg[3]), .A2(i_reg[10]), .A3(n175), .Z(N32) );
  nd02d1 U219 ( .A1(n172), .A2(n171), .ZN(n173) );
  xr03d1 U220 ( .A1(n172), .A2(i_reg[2]), .A3(n171), .Z(N31) );
  xr03d1 U221 ( .A1(i_reg[8]), .A2(i_reg[1]), .A3(n2), .Z(n1) );
  an02d1 U222 ( .A1(i_reg[0]), .A2(i_reg[7]), .Z(n2) );
  nr03d0 U223 ( .A1(n81), .A2(n131), .A3(n160), .ZN(n165) );
  an02d1 U224 ( .A1(i_reg[7]), .A2(i_reg[0]), .Z(n170) );
  cg01d1 U225 ( .A(i_reg[1]), .B(i_reg[8]), .CI(n170), .CO(n174) );
  xr02d1 U226 ( .A1(i_reg[0]), .A2(i_reg[7]), .Z(N29) );
  aor22d1 U227 ( .A1(i_reg[9]), .A2(n174), .B1(i_reg[2]), .B2(n173), .Z(n175)
         );
endmodule


module PCI_TOP ( pclk, pci_rst_n, pidsel, pgnt_n, pad_in, pad_out, pad_en, 
        ppar_in, ppar_out, ppar_en, pc_be_in, pc_be_out, pc_be_en, pframe_n_in, 
        pframe_n_out, pframe_n_en, ptrdy_n_in, ptrdy_n_out, ptrdy_n_en, 
        pirdy_n_in, pirdy_n_out, pirdy_n_en, pdevsel_n_in, pdevsel_n_out, 
        pdevsel_n_en, pstop_n_in, pstop_n_out, pstop_n_en, pperr_n_in, 
        pperr_n_out, pperr_n_en, pserr_n_in, pserr_n_out, pserr_n_en, preq_n, 
        pm66en, cmd_valid, cmd, cmd_in_valid, cmd_in, sys_clk, sys_rst_n, 
        test_mode, rfifo_pop, rfifo_empty, wfifo_push, wfifo_full, 
        pci_read_data, pci_write_data, test_si1, test_si2, test_si3, test_se, 
        test_so2, test_so3 );
  input [15:0] pad_in;
  output [15:0] pad_out;
  input [3:0] pc_be_in;
  output [3:0] pc_be_out;
  output [3:0] cmd;
  input [3:0] cmd_in;
  output [31:0] pci_read_data;
  input [31:0] pci_write_data;
  input pclk, pci_rst_n, pidsel, pgnt_n, ppar_in, pframe_n_in, ptrdy_n_in,
         pirdy_n_in, pdevsel_n_in, pstop_n_in, pperr_n_in, pserr_n_in, pm66en,
         cmd_in_valid, sys_clk, sys_rst_n, test_mode, rfifo_pop, wfifo_push,
         test_si1, test_si2, test_si3, test_se;
  output pad_en, ppar_out, ppar_en, pc_be_en, pframe_n_out, pframe_n_en,
         ptrdy_n_out, ptrdy_n_en, pirdy_n_out, pirdy_n_en, pdevsel_n_out,
         pdevsel_n_en, pstop_n_out, pstop_n_en, pperr_n_out, pperr_n_en,
         pserr_n_out, pserr_n_en, preq_n, cmd_valid, rfifo_empty, wfifo_full,
         test_so2, test_so3;
  wire   net_pci_read_push, net_pci_read_full, net_pci_write_pop,
         net_pci_write_empty, n3, n6, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40;
  wire   [31:0] net_pci_read_data;
  wire   [31:0] net_pci_write_data;

  PCI_CORE I_PCI_CORE ( .pclk(pclk), .pci_rst_n(pci_rst_n), .pidsel(pidsel), 
        .pgnt_n(pgnt_n), .pad_in(pad_in), .pad_out(pad_out), .pad_en(pad_en), 
        .ppar_in(ppar_in), .ppar_out(ppar_out), .ppar_en(ppar_en), .pc_be_in(
        pc_be_in), .pc_be_out(pc_be_out), .pc_be_en(pc_be_en), .pframe_n_in(
        pframe_n_in), .pframe_n_out(pframe_n_out), .pframe_n_en(pframe_n_en), 
        .ptrdy_n_in(ptrdy_n_in), .ptrdy_n_out(ptrdy_n_out), .ptrdy_n_en(
        ptrdy_n_en), .pirdy_n_in(pirdy_n_in), .pirdy_n_out(pirdy_n_out), 
        .pirdy_n_en(pirdy_n_en), .pdevsel_n_in(pdevsel_n_in), .pdevsel_n_out(
        pdevsel_n_out), .pdevsel_n_en(pdevsel_n_en), .pstop_n_in(pstop_n_in), 
        .pstop_n_out(pstop_n_out), .pstop_n_en(pstop_n_en), .pperr_n_in(
        pperr_n_in), .pperr_n_out(pperr_n_out), .pperr_n_en(pperr_n_en), 
        .pserr_n_in(pserr_n_in), .pserr_n_out(pserr_n_out), .pserr_n_en(
        pserr_n_en), .preq_n(preq_n), .pm66en(pm66en), .read_data(
        net_pci_read_data), .write_data(net_pci_write_data), .read_push(
        net_pci_read_push), .read_full(net_pci_read_full), .write_pop(
        net_pci_write_pop), .write_empty(net_pci_write_empty), .cmd_valid(
        cmd_valid), .cmd(cmd), .cmd_in_valid(cmd_in_valid), .cmd_in(cmd_in), 
        .test_se(test_se), .test_si1(test_si1), .test_si2(test_si2) );
  PCI_FIFO_0 I_PCI_READ_FIFO ( .fifo_clk_push(pclk), .fifo_clk_pop(sys_clk), 
        .fifo_rst_n(pci_rst_n), .test_mode(test_mode), .fifo_push_req_n(
        net_pci_read_push), .fifo_pop_req_n(rfifo_pop), .fifo_data_in(
        net_pci_read_data), .push_empty_fifo(SYNOPSYS_UNCONNECTED_21), 
        .push_ae_fifo(SYNOPSYS_UNCONNECTED_22), .push_hf_fifo(
        SYNOPSYS_UNCONNECTED_23), .push_af_fifo(SYNOPSYS_UNCONNECTED_24), 
        .push_full_fifo(net_pci_read_full), .push_error_fifo(
        SYNOPSYS_UNCONNECTED_25), .pop_empty_fifo(rfifo_empty), .pop_ae_fifo(
        SYNOPSYS_UNCONNECTED_26), .pop_hf_fifo(SYNOPSYS_UNCONNECTED_27), 
        .pop_af_fifo(SYNOPSYS_UNCONNECTED_28), .pop_full_fifo(
        SYNOPSYS_UNCONNECTED_29), .pop_error_fifo(SYNOPSYS_UNCONNECTED_30), 
        .data_out_fifo(pci_read_data), .test_si1(pc_be_en), .test_si2(test_si3), .test_se(test_se), .test_so1(n6), .test_so2(n3) );
  PCI_FIFO_1 I_PCI_WRITE_FIFO ( .fifo_clk_push(sys_clk), .fifo_clk_pop(pclk), 
        .fifo_rst_n(sys_rst_n), .test_mode(test_mode), .fifo_push_req_n(
        wfifo_push), .fifo_pop_req_n(net_pci_write_pop), .fifo_data_in(
        pci_write_data), .push_empty_fifo(SYNOPSYS_UNCONNECTED_31), 
        .push_ae_fifo(SYNOPSYS_UNCONNECTED_32), .push_hf_fifo(
        SYNOPSYS_UNCONNECTED_33), .push_af_fifo(SYNOPSYS_UNCONNECTED_34), 
        .push_full_fifo(wfifo_full), .push_error_fifo(SYNOPSYS_UNCONNECTED_35), 
        .pop_empty_fifo(net_pci_write_empty), .pop_ae_fifo(
        SYNOPSYS_UNCONNECTED_36), .pop_hf_fifo(SYNOPSYS_UNCONNECTED_37), 
        .pop_af_fifo(SYNOPSYS_UNCONNECTED_38), .pop_full_fifo(
        SYNOPSYS_UNCONNECTED_39), .pop_error_fifo(SYNOPSYS_UNCONNECTED_40), 
        .data_out_fifo(net_pci_write_data), .test_si1(n6), .test_si2(n3), 
        .test_se(test_se), .test_so1(test_so2), .test_so2(test_so3) );
endmodule


module ORCA_TOP ( sys_clk, sys_2x_clk, sdram_clk, scan_en, test_mode, 
        pci_rst_n, sdram_rst_n, sys_rst_n, sys_2x_rst_n, pclk, pidsel, pgnt_n, 
        pad_in, pad_out, pad_en, ppar_in, ppar_out, ppar_en, pc_be_in, 
        pc_be_out, pc_be_en, pframe_n_in, pframe_n_out, pframe_n_en, 
        ptrdy_n_in, ptrdy_n_out, ptrdy_n_en, pirdy_n_in, pirdy_n_out, 
        pirdy_n_en, pdevsel_n_in, pdevsel_n_out, pdevsel_n_en, pstop_n_in, 
        pstop_n_out, pstop_n_en, pperr_n_in, pperr_n_out, pperr_n_en, 
        pserr_n_in, pserr_n_out, pserr_n_en, preq_n, pm66en, sd_A, sd_CK, 
        sd_CKn, sd_LD, sd_RW, sd_BWS, sd_DQ_in, sd_DQ_out, sd_DQ_en );
  input [15:0] pad_in;
  output [15:0] pad_out;
  input [3:0] pc_be_in;
  output [3:0] pc_be_out;
  output [9:0] sd_A;
  output [1:0] sd_BWS;
  input [15:0] sd_DQ_in;
  output [15:0] sd_DQ_out;
  output [15:0] sd_DQ_en;
  input sys_clk, sys_2x_clk, sdram_clk, scan_en, test_mode, pci_rst_n,
         sdram_rst_n, sys_rst_n, sys_2x_rst_n, pclk, pidsel, pgnt_n, ppar_in,
         pframe_n_in, ptrdy_n_in, pirdy_n_in, pdevsel_n_in, pstop_n_in,
         pperr_n_in, pserr_n_in, pm66en;
  output pad_en, ppar_out, ppar_en, pc_be_en, pframe_n_out, pframe_n_en,
         ptrdy_n_out, ptrdy_n_en, pirdy_n_out, pirdy_n_en, pdevsel_n_out,
         pdevsel_n_en, pstop_n_out, pstop_n_en, pperr_n_out, pperr_n_en,
         pserr_n_out, pserr_n_en, preq_n, sd_CK, sd_CKn, sd_LD, sd_RW;
  wire   n18, n19, n20, n21, n22, n23, net_pci_parser_cmd_valid,
         net_parser_pci_cmd_valid, net_parser_fifo_read_pop,
         net_parser_fifo_read_empty, net_parser_fifo_write_push,
         net_parser_fifo_write_full, net_context_en, net_blender_clk_en,
         net_parser_sd_rfifo_pop, net_sd_rfifo_parser_empty,
         net_parser_sd_wfifo_push, net_sd_wfifo_parser_full,
         net_risc_sd_EndOfInstrn, net_risc_sd_Rd_Instr, net_risc_sd_OUT_VALID,
         net_risc_sd_STACK_FULL, net_blender_result_0__31_,
         net_blender_result_0__30_, net_blender_result_0__29_,
         net_blender_result_0__28_, net_blender_result_0__27_,
         net_blender_result_0__26_, net_blender_result_0__25_,
         net_blender_result_0__24_, net_blender_result_0__23_,
         net_blender_result_0__22_, net_blender_result_0__21_,
         net_blender_result_0__20_, net_blender_result_0__19_,
         net_blender_result_0__18_, net_blender_result_0__17_,
         net_blender_result_0__16_, net_blender_result_0__15_,
         net_blender_result_0__14_, net_blender_result_0__13_,
         net_blender_result_0__12_, net_blender_result_0__11_,
         net_blender_result_0__10_, net_blender_result_0__9_,
         net_blender_result_0__8_, net_blender_result_0__7_,
         net_blender_result_0__6_, net_blender_result_0__5_,
         net_blender_result_0__4_, net_blender_result_0__3_,
         net_blender_result_0__2_, net_blender_result_0__1_,
         net_blender_result_0__0_, n2, n5, n6, n7, n9, n11, n13, n14, n15, n17
;
  wire   [3:0] net_pci_parser_cmd;
  wire   [3:0] net_parser_pci_cmd;
  wire   [31:0] net_pci_sys_read_data;
  wire   [31:0] net_pci_wfifo_data;
  wire   [7:0] net_context_cmd;
  wire   [3:0] net_blender_op;
  wire   [7:0] net_parser_risc_Instrn_lo;
  wire   [31:0] net_risc_Xecutng_Instrn;
  wire   [1:0] net_pci_w_mux_select;
  wire   [1:0] net_sd_w_mux_select;
  wire   [31:0] net_pci_context_data;
  wire   [10:0] net_risc_sd_PSW;
  wire   [15:0] net_risc_RESULT_DATA;
  wire   [31:0] net_sd_sys_read_data;
  wire   [31:0] net_sd_wfifo_data;

  PCI_TOP I_PCI_TOP ( .pclk(pclk), .pci_rst_n(pci_rst_n), .pidsel(pidsel), 
        .pgnt_n(pgnt_n), .pad_in(pad_in), .pad_out(pad_out), .pad_en(pad_en), 
        .ppar_in(ppar_in), .ppar_out(ppar_out), .ppar_en(ppar_en), .pc_be_in(
        pc_be_in), .pc_be_out(pc_be_out), .pc_be_en(pc_be_en), .pframe_n_in(
        pframe_n_in), .pframe_n_out(pframe_n_out), .pframe_n_en(pframe_n_en), 
        .ptrdy_n_in(ptrdy_n_in), .ptrdy_n_out(ptrdy_n_out), .ptrdy_n_en(
        ptrdy_n_en), .pirdy_n_in(pirdy_n_in), .pirdy_n_out(pirdy_n_out), 
        .pirdy_n_en(pirdy_n_en), .pdevsel_n_in(pdevsel_n_in), .pdevsel_n_out(
        pdevsel_n_out), .pdevsel_n_en(pdevsel_n_en), .pstop_n_in(pstop_n_in), 
        .pstop_n_out(pstop_n_out), .pstop_n_en(pstop_n_en), .pperr_n_in(
        pperr_n_in), .pperr_n_out(pperr_n_out), .pperr_n_en(pperr_n_en), 
        .pserr_n_in(pserr_n_in), .pserr_n_out(pserr_n_out), .pserr_n_en(
        pserr_n_en), .preq_n(preq_n), .pm66en(pm66en), .cmd_valid(
        net_pci_parser_cmd_valid), .cmd(net_pci_parser_cmd), .cmd_in_valid(
        net_parser_pci_cmd_valid), .cmd_in(net_parser_pci_cmd), .sys_clk(
        sys_clk), .sys_rst_n(sys_rst_n), .test_mode(test_mode), .rfifo_pop(
        net_parser_fifo_read_pop), .rfifo_empty(net_parser_fifo_read_empty), 
        .wfifo_push(net_parser_fifo_write_push), .wfifo_full(
        net_parser_fifo_write_full), .pci_read_data(net_pci_sys_read_data), 
        .pci_write_data(net_pci_wfifo_data), .test_si1(n13), .test_si2(
        pad_in[2]), .test_si3(n6), .test_se(scan_en), .test_so2(n11), 
        .test_so3(n5) );
  PARSER I_PARSER ( .sys_clk(sys_clk), .pclk(pclk), .sys_rst_n(sys_rst_n), 
        .pcmd(net_pci_parser_cmd), .pcmd_valid(net_pci_parser_cmd_valid), 
        .pcmd_out(net_parser_pci_cmd), .pcmd_out_valid(
        net_parser_pci_cmd_valid), .blender_op(net_blender_op), 
        .blender_clk_en(net_blender_clk_en), .context_en(net_context_en), 
        .context_cmd(net_context_cmd), .fifo_read_pop(net_parser_fifo_read_pop), .fifo_read_empty(net_parser_fifo_read_empty), .fifo_write_push(
        net_parser_fifo_write_push), .fifo_write_full(
        net_parser_fifo_write_full), .risc_Instrn_lo(net_parser_risc_Instrn_lo), .risc_Xecutng_Instrn_lo(net_risc_Xecutng_Instrn[15:0]), .pci_w_mux_select(
        net_pci_w_mux_select), .sd_w_mux_select(net_sd_w_mux_select), 
        .parser_sd_rfifo_pop(net_parser_sd_rfifo_pop), .sd_rfifo_parser_empty(
        net_sd_rfifo_parser_empty), .parser_sd_wfifo_push(
        net_parser_sd_wfifo_push), .sd_wfifo_parser_full(
        net_sd_wfifo_parser_full), .test_se(scan_en), .test_si1(n7), 
        .test_si2(n14), .test_so2(n13), .test_so1(n6) );
  CONTEXT_MEM I_CONTEXT_MEM ( .sys_clk(sys_clk), .sys_rst_n(sys_rst_n), 
        .context_en(net_context_en), .cmd(net_context_cmd), .pci_data_in(
        net_pci_sys_read_data), .pci_context_data(net_pci_context_data) );
  RISC_CORE I_RISC_CORE ( .clk(sys_2x_clk), .reset_n(sys_2x_rst_n), .Instrn({
        net_pci_context_data[31:8], net_parser_risc_Instrn_lo}), 
        .Xecutng_Instrn(net_risc_Xecutng_Instrn), .EndOfInstrn(
        net_risc_sd_EndOfInstrn), .PSW(net_risc_sd_PSW), .Rd_Instr(
        net_risc_sd_Rd_Instr), .RESULT_DATA(net_risc_RESULT_DATA), .OUT_VALID(
        net_risc_sd_OUT_VALID), .STACK_FULL(net_risc_sd_STACK_FULL), 
        .test_si1(n9), .test_si2(pad_in[4]), .test_se(scan_en), .test_so2(n7)
         );
  BLENDER I_BLENDER_1 ( .clk(sys_clk), .reset_n(sys_rst_n), .clk_enable(
        net_blender_clk_en), .test_mode(test_mode), .operation(net_blender_op), 
        .op1(net_sd_sys_read_data), .op2(net_pci_context_data), .result({
        net_blender_result_0__31_, net_blender_result_0__30_, 
        net_blender_result_0__29_, net_blender_result_0__28_, 
        net_blender_result_0__27_, net_blender_result_0__26_, 
        net_blender_result_0__25_, net_blender_result_0__24_, 
        net_blender_result_0__23_, net_blender_result_0__22_, 
        net_blender_result_0__21_, net_blender_result_0__20_, 
        net_blender_result_0__19_, net_blender_result_0__18_, 
        net_blender_result_0__17_, net_blender_result_0__16_, 
        net_blender_result_0__15_, net_blender_result_0__14_, 
        net_blender_result_0__13_, net_blender_result_0__12_, 
        net_blender_result_0__11_, net_blender_result_0__10_, 
        net_blender_result_0__9_, net_blender_result_0__8_, 
        net_blender_result_0__7_, net_blender_result_0__6_, 
        net_blender_result_0__5_, net_blender_result_0__4_, 
        net_blender_result_0__3_, net_blender_result_0__2_, 
        net_blender_result_0__1_, net_blender_result_0__0_}), .test_se(scan_en), .test_si1(n17), .test_si2(pad_in[1]), .test_so2(n14), .test_so1(n15) );
  SDRAM_TOP I_SDRAM_TOP ( .sys_clk(sys_clk), .sdram_clk(sdram_clk), 
        .sys_rst_n(sys_rst_n), .sdram_rst_n(sdram_rst_n), .test_mode(test_mode), .risc_OUT_VALID(net_risc_sd_OUT_VALID), .risc_STACK_FULL(
        net_risc_sd_STACK_FULL), .risc_EndOfInstrn(net_risc_sd_EndOfInstrn), 
        .risc_PSW(net_risc_sd_PSW), .risc_Rd_Instr(net_risc_sd_Rd_Instr), 
        .sd_A({sd_A[9:6], n18, n19, n20, n21, n22, n23}), .sd_CK(sd_CK), 
        .sd_CKn(sd_CKn), .sd_LD(sd_LD), .sd_RW(sd_RW), .sd_BWS(sd_BWS), 
        .sd_DQ_in(sd_DQ_in), .sd_DQ_out(sd_DQ_out), .sd_DQ_en(sd_DQ_en), 
        .sd_sys_data_out(net_sd_sys_read_data), .sd_wfifo_data(
        net_sd_wfifo_data), .parser_sd_rfifo_pop(net_parser_sd_rfifo_pop), 
        .parser_sd_wfifo_push(net_parser_sd_wfifo_push), 
        .sd_rfifo_parser_empty(net_sd_rfifo_parser_empty), 
        .sd_wfifo_parser_full(net_sd_wfifo_parser_full), .test_si1(pad_in[0]), 
        .test_si2(n11), .test_si3(pad_in[3]), .test_si4(n5), .test_si5(
        pad_in[5]), .test_se(scan_en), .test_so1(n17), .test_so3(n9), 
        .test_so5(n2) );
  PCI_W_MUX I_PCI_W_MUX ( .blender_data({net_blender_result_0__31_, 
        net_blender_result_0__30_, net_blender_result_0__29_, 
        net_blender_result_0__28_, net_blender_result_0__27_, 
        net_blender_result_0__26_, net_blender_result_0__25_, 
        net_blender_result_0__24_, net_blender_result_0__23_, 
        net_blender_result_0__22_, net_blender_result_0__21_, 
        net_blender_result_0__20_, net_blender_result_0__19_, 
        net_blender_result_0__18_, net_blender_result_0__17_, 
        net_blender_result_0__16_, net_blender_result_0__15_, 
        net_blender_result_0__14_, net_blender_result_0__13_, 
        net_blender_result_0__12_, net_blender_result_0__11_, 
        net_blender_result_0__10_, net_blender_result_0__9_, 
        net_blender_result_0__8_, net_blender_result_0__7_, 
        net_blender_result_0__6_, net_blender_result_0__5_, 
        net_blender_result_0__4_, net_blender_result_0__3_, 
        net_blender_result_0__2_, net_blender_result_0__1_, 
        net_blender_result_0__0_}), .sdram_read_data(net_sd_sys_read_data), 
        .risc_result_data({net_risc_RESULT_DATA, 
        net_risc_Xecutng_Instrn[31:16]}), .pci_w_select(net_pci_w_mux_select), 
        .pci_wfifo_data(net_pci_wfifo_data) );
  SD_W_MUX I_SD_W_MUX ( .blender_data({net_blender_result_0__31_, 
        net_blender_result_0__30_, net_blender_result_0__29_, 
        net_blender_result_0__28_, net_blender_result_0__27_, 
        net_blender_result_0__26_, net_blender_result_0__25_, 
        net_blender_result_0__24_, net_blender_result_0__23_, 
        net_blender_result_0__22_, net_blender_result_0__21_, 
        net_blender_result_0__20_, net_blender_result_0__19_, 
        net_blender_result_0__18_, net_blender_result_0__17_, 
        net_blender_result_0__16_, net_blender_result_0__15_, 
        net_blender_result_0__14_, net_blender_result_0__13_, 
        net_blender_result_0__12_, net_blender_result_0__11_, 
        net_blender_result_0__10_, net_blender_result_0__9_, 
        net_blender_result_0__8_, net_blender_result_0__7_, 
        net_blender_result_0__6_, net_blender_result_0__5_, 
        net_blender_result_0__4_, net_blender_result_0__3_, 
        net_blender_result_0__2_, net_blender_result_0__1_, 
        net_blender_result_0__0_}), .pci_read_data(net_pci_context_data), 
        .risc_result_data({net_risc_RESULT_DATA, 
        net_risc_Xecutng_Instrn[31:16]}), .sd_w_select(net_sd_w_mux_select), 
        .sd_wfifo_data(net_sd_wfifo_data) );
  mx02d0 DFTC_U1 ( .I0(n18), .I1(n2), .S(scan_en), .Z(sd_A[5]) );
  mx02d0 DFTC_U2 ( .I0(n19), .I1(net_sd_sys_read_data[9]), .S(scan_en), .Z(
        sd_A[4]) );
  mx02d0 DFTC_U3 ( .I0(n20), .I1(net_risc_Xecutng_Instrn[2]), .S(scan_en), .Z(
        sd_A[3]) );
  mx02d0 DFTC_U4 ( .I0(n21), .I1(sd_BWS[1]), .S(scan_en), .Z(sd_A[2]) );
  mx02d0 DFTC_U5 ( .I0(n22), .I1(pad_out[2]), .S(scan_en), .Z(sd_A[1]) );
  mx02d0 DFTC_U6 ( .I0(n23), .I1(n15), .S(scan_en), .Z(sd_A[0]) );
endmodule

