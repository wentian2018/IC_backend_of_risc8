* File: rcx_out.net
* Created: Tue Mar 26 09:51:13 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:51:13 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt DFFDRX1  CK D Q QN RN VDD VSS
* 
XM76/X1 net0122 D VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM4/X1 MA MD net089 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM56/X1 MD ck2n net0116 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM52/X1 net0138 R VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM50/X1 MC MB net0138 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM48/X1 net0119 MA VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM49/X1 MB ck1n net0119 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM58/X1 SA SD net0132 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM72/X1 SB ck1n net0112 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM65/X1 SD ck2p net0129 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM64/X1 net0129 SC VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM69/X1 QN SC VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM66/X1 QN SA VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM63/X1 net0130 R VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM68/X1 Q SD VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM67/X1 Q SB VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM60/X1 net0131 SA VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM59/X1 net0132 R VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM62/X1 SC SB net0130 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM71/X1 SD ck2n net0110 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM70/X1 net0110 MC VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM61/X1 SB ck1p net0131 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM73/X1 net0112 MA VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM75/X1 MD ck2p net0120 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM9/X1 net089 R VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8801e-12 PD=2.23088e-05
XM74/X1 net0120 D VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM54/X1 net0116 MC VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM77/X1 MB ck1p net0122 VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XM5/X1 MA R VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=5.0305e-12 PD=1.68688e-05
XM57/X1 QN SA VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM55/X1 Q SB VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM53/X1 QN SC VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM51/X1 Q SD VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM44/X1 SB ck1n net0135 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM45/X1 SD ck2n net0133 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM42/X1 SA R VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM16/X1 MC R VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM39/X1 SA SB VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM33/X1 net0133 SA VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM32/X1 net0135 SC VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM38/X1 SC SD VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM36/X1 SC R VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM30/X1 SD ck2p net0111 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM29/X1 net0111 MC VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM26/X1 net0113 MA VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM22/X1 MD ck2p net0117 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM21/X1 net0117 MA VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM8/X1 MC MD VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM23/X1 SB ck1p net0113 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM14/X1 MB ck1p net0118 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM13/X1 net0118 MC VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM10/X1 MA MB VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM7/X1 MD ck2n net0121 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM6/X1 net0121 D VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM3/X1 net4 D VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XM0/X1 MB ck1n net4 VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XI4/XM1/X1 R RN VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XI4/XM0/X1 R RN VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XI3/XM1/X1 ck2n CK VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XI3/XM0/X1 ck2n CK VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XI1/XM1/X1 ck2p ck2n VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XI1/XM0/X1 ck2p ck2n VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XI0/XM1/X1 ck1p ck1n VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XI0/XM0/X1 ck1p ck1n VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
XI2/XM1/X1 ck1n CK VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9795e-12 PD=1.68288e-05
XI2/XM0/X1 ck1n CK VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8019e-12 PD=2.22688e-05
*
* 
* .include "rcx_out.net.DFFDRX1.pxi"
* BEGIN of "./rcx_out.net.DFFDRX1.pxi"
* File: rcx_out.net.DFFDRX1.pxi
* Created: Tue Mar 26 09:51:13 2019
* 

* END of "./rcx_out.net.DFFDRX1.pxi"
* 
*
.ends
*
*

