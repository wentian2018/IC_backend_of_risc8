# For SMIC 65LL/55LL Logic 1.2/2.5/3.3V Process
# Metal option: 1P9M_8Ic_1TMc_ALPA1
# 
# Reference technology documents:
#   1. Design Rule:       TD-LO55-DR-2002     rev. 5
#   2. SPICE Model:       TD-LO55-SP-2002     rev. 4
# 
# Copyright (c) 2016-2018 Cogenda Pte Ltd
# 
# All rights reserved
# 

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;
NAMESCASESENSITIVE ON ;
USEMINSPACING OBS OFF ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;

LAYER AA
  TYPE MASTERSLICE ;
END AA

LAYER GT
  TYPE MASTERSLICE ;
END GT

LAYER CT
  TYPE CUT ;
END CT

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.09 ;
  MINWIDTH 0.09 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.09 0.09
    WIDTH 1.001 0.09 0.16
    WIDTH 5.001 0.09 0.5
    WIDTH 12.001 0.09 0.5 ;
  AREA 0.027 ;
  MINENCLOSEDAREA 0.13 ;
  MAXWIDTH 12 ;
END M1

LAYER V1
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M2

LAYER V2
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0.005 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M3

LAYER V3
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0.005 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M4

LAYER V4
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0.005 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M5

LAYER V5
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0.005 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M6

LAYER V6
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0.005 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M7

LAYER V7
  TYPE CUT ;
  WIDTH 0.09 ;
  SPACING 0.13 ;
  SPACING 0.11 SAMENET ;
  ENCLOSURE BELOW 0.03 0.005 ;
  ENCLOSURE ABOVE 0.02 0.005 ;
  ARRAYSPACING CUTSPACING 0.11 ARRAYCUTS 3 SPACING 0.15 ;
END V7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  OFFSET 0.1 ;
  WIDTH 0.1 ;
  MINWIDTH 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.1 0.1
    WIDTH 1.001 0.1 0.16
    WIDTH 5.001 0.1 0.5
    WIDTH 12.001 0.1 0.5 ;
  AREA 0.035 ;
  MINENCLOSEDAREA 0.12 ;
  MAXWIDTH 12 ;
END M8

LAYER TV2
  TYPE CUT ;
  WIDTH 0.36 ;
  SPACING 0.34 ;
  ENCLOSURE BELOW 0.05 0.01 ;
  ENCLOSURE ABOVE 0.02 0.02 ;
  ARRAYSPACING CUTSPACING 0.34 ARRAYCUTS 2 SPACING 0.56 ;
END TV2

LAYER TM2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.8 ;
  OFFSET 0.4 ;
  WIDTH 0.4 ;
  MINWIDTH 0.4 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 2.001
    WIDTH 0 0.4 0.4
    WIDTH 2.001 0.4 0.5 ;
  AREA 0.4 ;
  MINENCLOSEDAREA 0.6 ;
  MAXWIDTH 20 ;
END TM2

LAYER RDV
  TYPE CUT ;
  WIDTH 3 ;
  SPACING 3 ;
  ENCLOSURE BELOW 1 1 ;
  ENCLOSURE ABOVE 1.5 1.5 ;
END RDV

LAYER RDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 6 ;
  WIDTH 3 ;
  MINWIDTH 3 ;
  SPACING 3 ;
  AREA 9 ;
END RDL

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP
MAXVIASTACK 4 ;

VIA via1_HV DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.045 0.075 0.045 ;
  LAYER M2 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_HV

VIA via1_VH DEFAULT
  LAYER M1 ;
  RECT -0.045 -0.075 0.045 0.075 ;
  LAYER M2 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_VH

VIA via1_HH DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.045 0.075 0.045 ;
  LAYER M2 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_HH

VIA via1_VV DEFAULT
  LAYER M1 ;
  RECT -0.045 -0.075 0.045 0.075 ;
  LAYER M2 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_VV

VIA via2_VH DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M3 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_VH

VIA via2_HV DEFAULT
  LAYER M2 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M3 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_HV

VIA via2_VV DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M3 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_VV

VIA via2_HH DEFAULT
  LAYER M2 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M3 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_HH

VIA via3_HV DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M4 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_HV

VIA via3_VH DEFAULT
  LAYER M3 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M4 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_VH

VIA via3_HH DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M4 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_HH

VIA via3_VV DEFAULT
  LAYER M3 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M4 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_VV

VIA via4_VH DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M5 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_VH

VIA via4_HV DEFAULT
  LAYER M4 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M5 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_HV

VIA via4_VV DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M5 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_VV

VIA via4_HH DEFAULT
  LAYER M4 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M5 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_HH

VIA via5_HV DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M6 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_HV

VIA via5_VH DEFAULT
  LAYER M5 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M6 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_VH

VIA via5_HH DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M6 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_HH

VIA via5_VV DEFAULT
  LAYER M5 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M6 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_VV

VIA via6_VH DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M7 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_VH

VIA via6_HV DEFAULT
  LAYER M6 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M7 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_HV

VIA via6_VV DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M7 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_VV

VIA via6_HH DEFAULT
  LAYER M6 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M7 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_HH

VIA via7_HV DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M8 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_HV

VIA via7_VH DEFAULT
  LAYER M7 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M8 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_VH

VIA via7_HH DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.05 0.075 0.05 ;
  LAYER M8 ;
  RECT -0.065 -0.05 0.065 0.05 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_HH

VIA via7_VV DEFAULT
  LAYER M7 ;
  RECT -0.05 -0.075 0.05 0.075 ;
  LAYER M8 ;
  RECT -0.05 -0.065 0.05 0.065 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_VV

VIA via8_VX DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.23 0.19 0.23 ;
  LAYER TM2 ;
  RECT -0.2 -0.2 0.2 0.2 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
END via8_VX

VIA via8_HX DEFAULT
  LAYER M8 ;
  RECT -0.23 -0.19 0.23 0.19 ;
  LAYER TM2 ;
  RECT -0.2 -0.2 0.2 0.2 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
END via8_HX

VIA via9_RDV DEFAULT
  LAYER TM2 ;
  RECT -2.5 -2.5 2.5 2.5 ;
  LAYER RDL ;
  RECT -3 -3 3 3 ;
  LAYER RDV ;
  RECT -1.5 -1.5 1.5 1.5 ;
END via9_RDV

VIA via1_HV_X2H DEFAULT
  LAYER M1 ;
  RECT -0.175 -0.045 0.175 0.045 ;
  LAYER M2 ;
  RECT -0.15 -0.065 0.15 0.065 ;
  LAYER V1 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via1_HV_X2H

VIA via1_HV_X2E DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.045 0.275 0.045 ;
  LAYER M2 ;
  RECT -0.05 -0.065 0.25 0.065 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via1_HV_X2E

VIA via1_HV_X2W DEFAULT
  LAYER M1 ;
  RECT -0.275 -0.045 0.075 0.045 ;
  LAYER M2 ;
  RECT -0.25 -0.065 0.05 0.065 ;
  LAYER V1 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_HV_X2W

VIA via1_HV_X2V DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.145 0.075 0.145 ;
  LAYER M2 ;
  RECT -0.05 -0.165 0.05 0.165 ;
  LAYER V1 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via1_HV_X2V

VIA via1_HV_X2S DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.245 0.075 0.045 ;
  LAYER M2 ;
  RECT -0.05 -0.265 0.05 0.065 ;
  LAYER V1 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_HV_X2S

VIA via1_HV_X2N DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.045 0.075 0.245 ;
  LAYER M2 ;
  RECT -0.05 -0.065 0.05 0.265 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via1_HV_X2N

VIA via1_HV_X3H DEFAULT
  LAYER M1 ;
  RECT -0.275 -0.045 0.275 0.045 ;
  LAYER M2 ;
  RECT -0.25 -0.065 0.25 0.065 ;
  LAYER V1 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via1_HV_X3H

VIA via1_HV_X3E DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.045 0.475 0.045 ;
  LAYER M2 ;
  RECT -0.05 -0.065 0.45 0.065 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via1_HV_X3E

VIA via1_HV_X3W DEFAULT
  LAYER M1 ;
  RECT -0.475 -0.045 0.075 0.045 ;
  LAYER M2 ;
  RECT -0.45 -0.065 0.05 0.065 ;
  LAYER V1 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_HV_X3W

VIA via1_HV_X3V DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.245 0.075 0.245 ;
  LAYER M2 ;
  RECT -0.05 -0.265 0.05 0.265 ;
  LAYER V1 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via1_HV_X3V

VIA via1_HV_X3S DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.445 0.075 0.045 ;
  LAYER M2 ;
  RECT -0.05 -0.465 0.05 0.065 ;
  LAYER V1 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via1_HV_X3S

VIA via1_HV_X3N DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.045 0.075 0.445 ;
  LAYER M2 ;
  RECT -0.05 -0.065 0.05 0.465 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via1_HV_X3N

VIA via1_HV_X4H DEFAULT
  LAYER M1 ;
  RECT -0.175 -0.145 0.175 0.145 ;
  LAYER M2 ;
  RECT -0.15 -0.165 0.15 0.165 ;
  LAYER V1 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via1_HV_X4H

VIA via1_HV_X4E DEFAULT
  LAYER M1 ;
  RECT -0.075 -0.145 0.275 0.145 ;
  LAYER M2 ;
  RECT -0.05 -0.165 0.25 0.165 ;
  LAYER V1 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via1_HV_X4E

VIA via1_HV_X4W DEFAULT
  LAYER M1 ;
  RECT -0.275 -0.145 0.075 0.145 ;
  LAYER M2 ;
  RECT -0.25 -0.165 0.05 0.165 ;
  LAYER V1 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via1_HV_X4W

VIA via1_HV_X4S DEFAULT
  LAYER M1 ;
  RECT -0.175 -0.245 0.175 0.045 ;
  LAYER M2 ;
  RECT -0.15 -0.265 0.15 0.065 ;
  LAYER V1 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via1_HV_X4S

VIA via1_HV_X4N DEFAULT
  LAYER M1 ;
  RECT -0.175 -0.045 0.175 0.245 ;
  LAYER M2 ;
  RECT -0.15 -0.065 0.15 0.265 ;
  LAYER V1 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via1_HV_X4N

VIA via2_VH_X2H DEFAULT
  LAYER M2 ;
  RECT -0.15 -0.075 0.15 0.075 ;
  LAYER M3 ;
  RECT -0.165 -0.05 0.165 0.05 ;
  LAYER V2 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via2_VH_X2H

VIA via2_VH_X2E DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.075 0.25 0.075 ;
  LAYER M3 ;
  RECT -0.065 -0.05 0.265 0.05 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via2_VH_X2E

VIA via2_VH_X2W DEFAULT
  LAYER M2 ;
  RECT -0.25 -0.075 0.05 0.075 ;
  LAYER M3 ;
  RECT -0.265 -0.05 0.065 0.05 ;
  LAYER V2 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_VH_X2W

VIA via2_VH_X2V DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.175 0.05 0.175 ;
  LAYER M3 ;
  RECT -0.065 -0.15 0.065 0.15 ;
  LAYER V2 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via2_VH_X2V

VIA via2_VH_X2S DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.275 0.05 0.075 ;
  LAYER M3 ;
  RECT -0.065 -0.25 0.065 0.05 ;
  LAYER V2 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_VH_X2S

VIA via2_VH_X2N DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.075 0.05 0.275 ;
  LAYER M3 ;
  RECT -0.065 -0.05 0.065 0.25 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via2_VH_X2N

VIA via2_VH_X3H DEFAULT
  LAYER M2 ;
  RECT -0.25 -0.075 0.25 0.075 ;
  LAYER M3 ;
  RECT -0.265 -0.05 0.265 0.05 ;
  LAYER V2 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via2_VH_X3H

VIA via2_VH_X3E DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.075 0.45 0.075 ;
  LAYER M3 ;
  RECT -0.065 -0.05 0.465 0.05 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via2_VH_X3E

VIA via2_VH_X3W DEFAULT
  LAYER M2 ;
  RECT -0.45 -0.075 0.05 0.075 ;
  LAYER M3 ;
  RECT -0.465 -0.05 0.065 0.05 ;
  LAYER V2 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_VH_X3W

VIA via2_VH_X3V DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.275 0.05 0.275 ;
  LAYER M3 ;
  RECT -0.065 -0.25 0.065 0.25 ;
  LAYER V2 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via2_VH_X3V

VIA via2_VH_X3S DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.475 0.05 0.075 ;
  LAYER M3 ;
  RECT -0.065 -0.45 0.065 0.05 ;
  LAYER V2 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via2_VH_X3S

VIA via2_VH_X3N DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.075 0.05 0.475 ;
  LAYER M3 ;
  RECT -0.065 -0.05 0.065 0.45 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via2_VH_X3N

VIA via2_VH_X4H DEFAULT
  LAYER M2 ;
  RECT -0.15 -0.175 0.15 0.175 ;
  LAYER M3 ;
  RECT -0.165 -0.15 0.165 0.15 ;
  LAYER V2 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via2_VH_X4H

VIA via2_VH_X4E DEFAULT
  LAYER M2 ;
  RECT -0.05 -0.175 0.25 0.175 ;
  LAYER M3 ;
  RECT -0.065 -0.15 0.265 0.15 ;
  LAYER V2 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via2_VH_X4E

VIA via2_VH_X4W DEFAULT
  LAYER M2 ;
  RECT -0.25 -0.175 0.05 0.175 ;
  LAYER M3 ;
  RECT -0.265 -0.15 0.065 0.15 ;
  LAYER V2 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via2_VH_X4W

VIA via2_VH_X4S DEFAULT
  LAYER M2 ;
  RECT -0.15 -0.275 0.15 0.075 ;
  LAYER M3 ;
  RECT -0.165 -0.25 0.165 0.05 ;
  LAYER V2 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via2_VH_X4S

VIA via2_VH_X4N DEFAULT
  LAYER M2 ;
  RECT -0.15 -0.075 0.15 0.275 ;
  LAYER M3 ;
  RECT -0.165 -0.05 0.165 0.25 ;
  LAYER V2 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via2_VH_X4N

VIA via3_HV_X2H DEFAULT
  LAYER M3 ;
  RECT -0.175 -0.05 0.175 0.05 ;
  LAYER M4 ;
  RECT -0.15 -0.065 0.15 0.065 ;
  LAYER V3 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via3_HV_X2H

VIA via3_HV_X2E DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.05 0.275 0.05 ;
  LAYER M4 ;
  RECT -0.05 -0.065 0.25 0.065 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via3_HV_X2E

VIA via3_HV_X2W DEFAULT
  LAYER M3 ;
  RECT -0.275 -0.05 0.075 0.05 ;
  LAYER M4 ;
  RECT -0.25 -0.065 0.05 0.065 ;
  LAYER V3 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_HV_X2W

VIA via3_HV_X2V DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.15 0.075 0.15 ;
  LAYER M4 ;
  RECT -0.05 -0.165 0.05 0.165 ;
  LAYER V3 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via3_HV_X2V

VIA via3_HV_X2S DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.25 0.075 0.05 ;
  LAYER M4 ;
  RECT -0.05 -0.265 0.05 0.065 ;
  LAYER V3 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_HV_X2S

VIA via3_HV_X2N DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.05 0.075 0.25 ;
  LAYER M4 ;
  RECT -0.05 -0.065 0.05 0.265 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via3_HV_X2N

VIA via3_HV_X3H DEFAULT
  LAYER M3 ;
  RECT -0.275 -0.05 0.275 0.05 ;
  LAYER M4 ;
  RECT -0.25 -0.065 0.25 0.065 ;
  LAYER V3 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via3_HV_X3H

VIA via3_HV_X3E DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.05 0.475 0.05 ;
  LAYER M4 ;
  RECT -0.05 -0.065 0.45 0.065 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via3_HV_X3E

VIA via3_HV_X3W DEFAULT
  LAYER M3 ;
  RECT -0.475 -0.05 0.075 0.05 ;
  LAYER M4 ;
  RECT -0.45 -0.065 0.05 0.065 ;
  LAYER V3 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_HV_X3W

VIA via3_HV_X3V DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.25 0.075 0.25 ;
  LAYER M4 ;
  RECT -0.05 -0.265 0.05 0.265 ;
  LAYER V3 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via3_HV_X3V

VIA via3_HV_X3S DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.45 0.075 0.05 ;
  LAYER M4 ;
  RECT -0.05 -0.465 0.05 0.065 ;
  LAYER V3 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via3_HV_X3S

VIA via3_HV_X3N DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.05 0.075 0.45 ;
  LAYER M4 ;
  RECT -0.05 -0.065 0.05 0.465 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via3_HV_X3N

VIA via3_HV_X4H DEFAULT
  LAYER M3 ;
  RECT -0.175 -0.15 0.175 0.15 ;
  LAYER M4 ;
  RECT -0.15 -0.165 0.15 0.165 ;
  LAYER V3 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via3_HV_X4H

VIA via3_HV_X4E DEFAULT
  LAYER M3 ;
  RECT -0.075 -0.15 0.275 0.15 ;
  LAYER M4 ;
  RECT -0.05 -0.165 0.25 0.165 ;
  LAYER V3 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via3_HV_X4E

VIA via3_HV_X4W DEFAULT
  LAYER M3 ;
  RECT -0.275 -0.15 0.075 0.15 ;
  LAYER M4 ;
  RECT -0.25 -0.165 0.05 0.165 ;
  LAYER V3 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via3_HV_X4W

VIA via3_HV_X4S DEFAULT
  LAYER M3 ;
  RECT -0.175 -0.25 0.175 0.05 ;
  LAYER M4 ;
  RECT -0.15 -0.265 0.15 0.065 ;
  LAYER V3 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via3_HV_X4S

VIA via3_HV_X4N DEFAULT
  LAYER M3 ;
  RECT -0.175 -0.05 0.175 0.25 ;
  LAYER M4 ;
  RECT -0.15 -0.065 0.15 0.265 ;
  LAYER V3 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via3_HV_X4N

VIA via4_VH_X2H DEFAULT
  LAYER M4 ;
  RECT -0.15 -0.075 0.15 0.075 ;
  LAYER M5 ;
  RECT -0.165 -0.05 0.165 0.05 ;
  LAYER V4 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via4_VH_X2H

VIA via4_VH_X2E DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.075 0.25 0.075 ;
  LAYER M5 ;
  RECT -0.065 -0.05 0.265 0.05 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via4_VH_X2E

VIA via4_VH_X2W DEFAULT
  LAYER M4 ;
  RECT -0.25 -0.075 0.05 0.075 ;
  LAYER M5 ;
  RECT -0.265 -0.05 0.065 0.05 ;
  LAYER V4 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_VH_X2W

VIA via4_VH_X2V DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.175 0.05 0.175 ;
  LAYER M5 ;
  RECT -0.065 -0.15 0.065 0.15 ;
  LAYER V4 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via4_VH_X2V

VIA via4_VH_X2S DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.275 0.05 0.075 ;
  LAYER M5 ;
  RECT -0.065 -0.25 0.065 0.05 ;
  LAYER V4 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_VH_X2S

VIA via4_VH_X2N DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.075 0.05 0.275 ;
  LAYER M5 ;
  RECT -0.065 -0.05 0.065 0.25 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via4_VH_X2N

VIA via4_VH_X3H DEFAULT
  LAYER M4 ;
  RECT -0.25 -0.075 0.25 0.075 ;
  LAYER M5 ;
  RECT -0.265 -0.05 0.265 0.05 ;
  LAYER V4 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via4_VH_X3H

VIA via4_VH_X3E DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.075 0.45 0.075 ;
  LAYER M5 ;
  RECT -0.065 -0.05 0.465 0.05 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via4_VH_X3E

VIA via4_VH_X3W DEFAULT
  LAYER M4 ;
  RECT -0.45 -0.075 0.05 0.075 ;
  LAYER M5 ;
  RECT -0.465 -0.05 0.065 0.05 ;
  LAYER V4 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_VH_X3W

VIA via4_VH_X3V DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.275 0.05 0.275 ;
  LAYER M5 ;
  RECT -0.065 -0.25 0.065 0.25 ;
  LAYER V4 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via4_VH_X3V

VIA via4_VH_X3S DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.475 0.05 0.075 ;
  LAYER M5 ;
  RECT -0.065 -0.45 0.065 0.05 ;
  LAYER V4 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via4_VH_X3S

VIA via4_VH_X3N DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.075 0.05 0.475 ;
  LAYER M5 ;
  RECT -0.065 -0.05 0.065 0.45 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via4_VH_X3N

VIA via4_VH_X4H DEFAULT
  LAYER M4 ;
  RECT -0.15 -0.175 0.15 0.175 ;
  LAYER M5 ;
  RECT -0.165 -0.15 0.165 0.15 ;
  LAYER V4 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via4_VH_X4H

VIA via4_VH_X4E DEFAULT
  LAYER M4 ;
  RECT -0.05 -0.175 0.25 0.175 ;
  LAYER M5 ;
  RECT -0.065 -0.15 0.265 0.15 ;
  LAYER V4 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via4_VH_X4E

VIA via4_VH_X4W DEFAULT
  LAYER M4 ;
  RECT -0.25 -0.175 0.05 0.175 ;
  LAYER M5 ;
  RECT -0.265 -0.15 0.065 0.15 ;
  LAYER V4 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via4_VH_X4W

VIA via4_VH_X4S DEFAULT
  LAYER M4 ;
  RECT -0.15 -0.275 0.15 0.075 ;
  LAYER M5 ;
  RECT -0.165 -0.25 0.165 0.05 ;
  LAYER V4 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via4_VH_X4S

VIA via4_VH_X4N DEFAULT
  LAYER M4 ;
  RECT -0.15 -0.075 0.15 0.275 ;
  LAYER M5 ;
  RECT -0.165 -0.05 0.165 0.25 ;
  LAYER V4 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via4_VH_X4N

VIA via5_HV_X2H DEFAULT
  LAYER M5 ;
  RECT -0.175 -0.05 0.175 0.05 ;
  LAYER M6 ;
  RECT -0.15 -0.065 0.15 0.065 ;
  LAYER V5 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via5_HV_X2H

VIA via5_HV_X2E DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.05 0.275 0.05 ;
  LAYER M6 ;
  RECT -0.05 -0.065 0.25 0.065 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via5_HV_X2E

VIA via5_HV_X2W DEFAULT
  LAYER M5 ;
  RECT -0.275 -0.05 0.075 0.05 ;
  LAYER M6 ;
  RECT -0.25 -0.065 0.05 0.065 ;
  LAYER V5 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_HV_X2W

VIA via5_HV_X2V DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.15 0.075 0.15 ;
  LAYER M6 ;
  RECT -0.05 -0.165 0.05 0.165 ;
  LAYER V5 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via5_HV_X2V

VIA via5_HV_X2S DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.25 0.075 0.05 ;
  LAYER M6 ;
  RECT -0.05 -0.265 0.05 0.065 ;
  LAYER V5 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_HV_X2S

VIA via5_HV_X2N DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.05 0.075 0.25 ;
  LAYER M6 ;
  RECT -0.05 -0.065 0.05 0.265 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via5_HV_X2N

VIA via5_HV_X3H DEFAULT
  LAYER M5 ;
  RECT -0.275 -0.05 0.275 0.05 ;
  LAYER M6 ;
  RECT -0.25 -0.065 0.25 0.065 ;
  LAYER V5 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via5_HV_X3H

VIA via5_HV_X3E DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.05 0.475 0.05 ;
  LAYER M6 ;
  RECT -0.05 -0.065 0.45 0.065 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via5_HV_X3E

VIA via5_HV_X3W DEFAULT
  LAYER M5 ;
  RECT -0.475 -0.05 0.075 0.05 ;
  LAYER M6 ;
  RECT -0.45 -0.065 0.05 0.065 ;
  LAYER V5 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_HV_X3W

VIA via5_HV_X3V DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.25 0.075 0.25 ;
  LAYER M6 ;
  RECT -0.05 -0.265 0.05 0.265 ;
  LAYER V5 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via5_HV_X3V

VIA via5_HV_X3S DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.45 0.075 0.05 ;
  LAYER M6 ;
  RECT -0.05 -0.465 0.05 0.065 ;
  LAYER V5 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via5_HV_X3S

VIA via5_HV_X3N DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.05 0.075 0.45 ;
  LAYER M6 ;
  RECT -0.05 -0.065 0.05 0.465 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via5_HV_X3N

VIA via5_HV_X4H DEFAULT
  LAYER M5 ;
  RECT -0.175 -0.15 0.175 0.15 ;
  LAYER M6 ;
  RECT -0.15 -0.165 0.15 0.165 ;
  LAYER V5 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via5_HV_X4H

VIA via5_HV_X4E DEFAULT
  LAYER M5 ;
  RECT -0.075 -0.15 0.275 0.15 ;
  LAYER M6 ;
  RECT -0.05 -0.165 0.25 0.165 ;
  LAYER V5 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via5_HV_X4E

VIA via5_HV_X4W DEFAULT
  LAYER M5 ;
  RECT -0.275 -0.15 0.075 0.15 ;
  LAYER M6 ;
  RECT -0.25 -0.165 0.05 0.165 ;
  LAYER V5 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via5_HV_X4W

VIA via5_HV_X4S DEFAULT
  LAYER M5 ;
  RECT -0.175 -0.25 0.175 0.05 ;
  LAYER M6 ;
  RECT -0.15 -0.265 0.15 0.065 ;
  LAYER V5 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via5_HV_X4S

VIA via5_HV_X4N DEFAULT
  LAYER M5 ;
  RECT -0.175 -0.05 0.175 0.25 ;
  LAYER M6 ;
  RECT -0.15 -0.065 0.15 0.265 ;
  LAYER V5 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via5_HV_X4N

VIA via6_VH_X2H DEFAULT
  LAYER M6 ;
  RECT -0.15 -0.075 0.15 0.075 ;
  LAYER M7 ;
  RECT -0.165 -0.05 0.165 0.05 ;
  LAYER V6 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via6_VH_X2H

VIA via6_VH_X2E DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.075 0.25 0.075 ;
  LAYER M7 ;
  RECT -0.065 -0.05 0.265 0.05 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via6_VH_X2E

VIA via6_VH_X2W DEFAULT
  LAYER M6 ;
  RECT -0.25 -0.075 0.05 0.075 ;
  LAYER M7 ;
  RECT -0.265 -0.05 0.065 0.05 ;
  LAYER V6 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_VH_X2W

VIA via6_VH_X2V DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.175 0.05 0.175 ;
  LAYER M7 ;
  RECT -0.065 -0.15 0.065 0.15 ;
  LAYER V6 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via6_VH_X2V

VIA via6_VH_X2S DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.275 0.05 0.075 ;
  LAYER M7 ;
  RECT -0.065 -0.25 0.065 0.05 ;
  LAYER V6 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_VH_X2S

VIA via6_VH_X2N DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.075 0.05 0.275 ;
  LAYER M7 ;
  RECT -0.065 -0.05 0.065 0.25 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via6_VH_X2N

VIA via6_VH_X3H DEFAULT
  LAYER M6 ;
  RECT -0.25 -0.075 0.25 0.075 ;
  LAYER M7 ;
  RECT -0.265 -0.05 0.265 0.05 ;
  LAYER V6 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via6_VH_X3H

VIA via6_VH_X3E DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.075 0.45 0.075 ;
  LAYER M7 ;
  RECT -0.065 -0.05 0.465 0.05 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via6_VH_X3E

VIA via6_VH_X3W DEFAULT
  LAYER M6 ;
  RECT -0.45 -0.075 0.05 0.075 ;
  LAYER M7 ;
  RECT -0.465 -0.05 0.065 0.05 ;
  LAYER V6 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_VH_X3W

VIA via6_VH_X3V DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.275 0.05 0.275 ;
  LAYER M7 ;
  RECT -0.065 -0.25 0.065 0.25 ;
  LAYER V6 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via6_VH_X3V

VIA via6_VH_X3S DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.475 0.05 0.075 ;
  LAYER M7 ;
  RECT -0.065 -0.45 0.065 0.05 ;
  LAYER V6 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via6_VH_X3S

VIA via6_VH_X3N DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.075 0.05 0.475 ;
  LAYER M7 ;
  RECT -0.065 -0.05 0.065 0.45 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via6_VH_X3N

VIA via6_VH_X4H DEFAULT
  LAYER M6 ;
  RECT -0.15 -0.175 0.15 0.175 ;
  LAYER M7 ;
  RECT -0.165 -0.15 0.165 0.15 ;
  LAYER V6 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via6_VH_X4H

VIA via6_VH_X4E DEFAULT
  LAYER M6 ;
  RECT -0.05 -0.175 0.25 0.175 ;
  LAYER M7 ;
  RECT -0.065 -0.15 0.265 0.15 ;
  LAYER V6 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via6_VH_X4E

VIA via6_VH_X4W DEFAULT
  LAYER M6 ;
  RECT -0.25 -0.175 0.05 0.175 ;
  LAYER M7 ;
  RECT -0.265 -0.15 0.065 0.15 ;
  LAYER V6 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via6_VH_X4W

VIA via6_VH_X4S DEFAULT
  LAYER M6 ;
  RECT -0.15 -0.275 0.15 0.075 ;
  LAYER M7 ;
  RECT -0.165 -0.25 0.165 0.05 ;
  LAYER V6 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via6_VH_X4S

VIA via6_VH_X4N DEFAULT
  LAYER M6 ;
  RECT -0.15 -0.075 0.15 0.275 ;
  LAYER M7 ;
  RECT -0.165 -0.05 0.165 0.25 ;
  LAYER V6 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via6_VH_X4N

VIA via7_HV_X2H DEFAULT
  LAYER M7 ;
  RECT -0.175 -0.05 0.175 0.05 ;
  LAYER M8 ;
  RECT -0.15 -0.065 0.15 0.065 ;
  LAYER V7 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via7_HV_X2H

VIA via7_HV_X2E DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.05 0.275 0.05 ;
  LAYER M8 ;
  RECT -0.05 -0.065 0.25 0.065 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via7_HV_X2E

VIA via7_HV_X2W DEFAULT
  LAYER M7 ;
  RECT -0.275 -0.05 0.075 0.05 ;
  LAYER M8 ;
  RECT -0.25 -0.065 0.05 0.065 ;
  LAYER V7 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_HV_X2W

VIA via7_HV_X2V DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.15 0.075 0.15 ;
  LAYER M8 ;
  RECT -0.05 -0.165 0.05 0.165 ;
  LAYER V7 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via7_HV_X2V

VIA via7_HV_X2S DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.25 0.075 0.05 ;
  LAYER M8 ;
  RECT -0.05 -0.265 0.05 0.065 ;
  LAYER V7 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_HV_X2S

VIA via7_HV_X2N DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.05 0.075 0.25 ;
  LAYER M8 ;
  RECT -0.05 -0.065 0.05 0.265 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via7_HV_X2N

VIA via7_HV_X3H DEFAULT
  LAYER M7 ;
  RECT -0.275 -0.05 0.275 0.05 ;
  LAYER M8 ;
  RECT -0.25 -0.065 0.25 0.065 ;
  LAYER V7 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
END via7_HV_X3H

VIA via7_HV_X3E DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.05 0.475 0.05 ;
  LAYER M8 ;
  RECT -0.05 -0.065 0.45 0.065 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT 0.155 -0.045 0.245 0.045 ;
  RECT 0.355 -0.045 0.445 0.045 ;
END via7_HV_X3E

VIA via7_HV_X3W DEFAULT
  LAYER M7 ;
  RECT -0.475 -0.05 0.075 0.05 ;
  LAYER M8 ;
  RECT -0.45 -0.065 0.05 0.065 ;
  LAYER V7 ;
  RECT -0.445 -0.045 -0.355 0.045 ;
  RECT -0.245 -0.045 -0.155 0.045 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_HV_X3W

VIA via7_HV_X3V DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.25 0.075 0.25 ;
  LAYER M8 ;
  RECT -0.05 -0.265 0.05 0.265 ;
  LAYER V7 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
END via7_HV_X3V

VIA via7_HV_X3S DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.45 0.075 0.05 ;
  LAYER M8 ;
  RECT -0.05 -0.465 0.05 0.065 ;
  LAYER V7 ;
  RECT -0.045 -0.445 0.045 -0.355 ;
  RECT -0.045 -0.245 0.045 -0.155 ;
  RECT -0.045 -0.045 0.045 0.045 ;
END via7_HV_X3S

VIA via7_HV_X3N DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.05 0.075 0.45 ;
  LAYER M8 ;
  RECT -0.05 -0.065 0.05 0.465 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  RECT -0.045 0.155 0.045 0.245 ;
  RECT -0.045 0.355 0.045 0.445 ;
END via7_HV_X3N

VIA via7_HV_X4H DEFAULT
  LAYER M7 ;
  RECT -0.175 -0.15 0.175 0.15 ;
  LAYER M8 ;
  RECT -0.15 -0.165 0.15 0.165 ;
  LAYER V7 ;
  RECT -0.145 -0.145 -0.055 -0.055 ;
  RECT -0.145 0.055 -0.055 0.145 ;
  RECT 0.055 -0.145 0.145 -0.055 ;
  RECT 0.055 0.055 0.145 0.145 ;
END via7_HV_X4H

VIA via7_HV_X4E DEFAULT
  LAYER M7 ;
  RECT -0.075 -0.15 0.275 0.15 ;
  LAYER M8 ;
  RECT -0.05 -0.165 0.25 0.165 ;
  LAYER V7 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
  RECT 0.155 -0.145 0.245 -0.055 ;
  RECT 0.155 0.055 0.245 0.145 ;
END via7_HV_X4E

VIA via7_HV_X4W DEFAULT
  LAYER M7 ;
  RECT -0.275 -0.15 0.075 0.15 ;
  LAYER M8 ;
  RECT -0.25 -0.165 0.05 0.165 ;
  LAYER V7 ;
  RECT -0.245 -0.145 -0.155 -0.055 ;
  RECT -0.245 0.055 -0.155 0.145 ;
  RECT -0.045 -0.145 0.045 -0.055 ;
  RECT -0.045 0.055 0.045 0.145 ;
END via7_HV_X4W

VIA via7_HV_X4S DEFAULT
  LAYER M7 ;
  RECT -0.175 -0.25 0.175 0.05 ;
  LAYER M8 ;
  RECT -0.15 -0.265 0.15 0.065 ;
  LAYER V7 ;
  RECT -0.145 -0.245 -0.055 -0.155 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT 0.055 -0.245 0.145 -0.155 ;
  RECT 0.055 -0.045 0.145 0.045 ;
END via7_HV_X4S

VIA via7_HV_X4N DEFAULT
  LAYER M7 ;
  RECT -0.175 -0.05 0.175 0.25 ;
  LAYER M8 ;
  RECT -0.15 -0.065 0.15 0.265 ;
  LAYER V7 ;
  RECT -0.145 -0.045 -0.055 0.045 ;
  RECT -0.145 0.155 -0.055 0.245 ;
  RECT 0.055 -0.045 0.145 0.045 ;
  RECT 0.055 0.155 0.145 0.245 ;
END via7_HV_X4N

VIA via8_VX_X2H DEFAULT
  LAYER M8 ;
  RECT -0.54 -0.23 0.54 0.23 ;
  LAYER TM2 ;
  RECT -0.55 -0.2 0.55 0.2 ;
  LAYER TV2 ;
  RECT -0.53 -0.18 -0.17 0.18 ;
  RECT 0.17 -0.18 0.53 0.18 ;
END via8_VX_X2H

VIA via8_VX_X2E DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.23 0.89 0.23 ;
  LAYER TM2 ;
  RECT -0.2 -0.2 0.9 0.2 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  RECT 0.52 -0.18 0.88 0.18 ;
END via8_VX_X2E

VIA via8_VX_X2W DEFAULT
  LAYER M8 ;
  RECT -0.89 -0.23 0.19 0.23 ;
  LAYER TM2 ;
  RECT -0.9 -0.2 0.2 0.2 ;
  LAYER TV2 ;
  RECT -0.88 -0.18 -0.52 0.18 ;
  RECT -0.18 -0.18 0.18 0.18 ;
END via8_VX_X2W

VIA via8_VX_X2V DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.58 0.19 0.58 ;
  LAYER TM2 ;
  RECT -0.2 -0.55 0.2 0.55 ;
  LAYER TV2 ;
  RECT -0.18 -0.53 0.18 -0.17 ;
  RECT -0.18 0.17 0.18 0.53 ;
END via8_VX_X2V

VIA via8_VX_X2S DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.93 0.19 0.23 ;
  LAYER TM2 ;
  RECT -0.2 -0.9 0.2 0.2 ;
  LAYER TV2 ;
  RECT -0.18 -0.88 0.18 -0.52 ;
  RECT -0.18 -0.18 0.18 0.18 ;
END via8_VX_X2S

VIA via8_VX_X2N DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.23 0.19 0.93 ;
  LAYER TM2 ;
  RECT -0.2 -0.2 0.2 0.9 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  RECT -0.18 0.52 0.18 0.88 ;
END via8_VX_X2N

VIA via8_VX_X3H DEFAULT
  LAYER M8 ;
  RECT -0.89 -0.23 0.89 0.23 ;
  LAYER TM2 ;
  RECT -0.9 -0.2 0.9 0.2 ;
  LAYER TV2 ;
  RECT -0.88 -0.18 -0.52 0.18 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  RECT 0.52 -0.18 0.88 0.18 ;
END via8_VX_X3H

VIA via8_VX_X3E DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.23 1.59 0.23 ;
  LAYER TM2 ;
  RECT -0.2 -0.2 1.6 0.2 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  RECT 0.52 -0.18 0.88 0.18 ;
  RECT 1.22 -0.18 1.58 0.18 ;
END via8_VX_X3E

VIA via8_VX_X3W DEFAULT
  LAYER M8 ;
  RECT -1.59 -0.23 0.19 0.23 ;
  LAYER TM2 ;
  RECT -1.6 -0.2 0.2 0.2 ;
  LAYER TV2 ;
  RECT -1.58 -0.18 -1.22 0.18 ;
  RECT -0.88 -0.18 -0.52 0.18 ;
  RECT -0.18 -0.18 0.18 0.18 ;
END via8_VX_X3W

VIA via8_VX_X3V DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.93 0.19 0.93 ;
  LAYER TM2 ;
  RECT -0.2 -0.9 0.2 0.9 ;
  LAYER TV2 ;
  RECT -0.18 -0.88 0.18 -0.52 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  RECT -0.18 0.52 0.18 0.88 ;
END via8_VX_X3V

VIA via8_VX_X3S DEFAULT
  LAYER M8 ;
  RECT -0.19 -1.63 0.19 0.23 ;
  LAYER TM2 ;
  RECT -0.2 -1.6 0.2 0.2 ;
  LAYER TV2 ;
  RECT -0.18 -1.58 0.18 -1.22 ;
  RECT -0.18 -0.88 0.18 -0.52 ;
  RECT -0.18 -0.18 0.18 0.18 ;
END via8_VX_X3S

VIA via8_VX_X3N DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.23 0.19 1.63 ;
  LAYER TM2 ;
  RECT -0.2 -0.2 0.2 1.6 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  RECT -0.18 0.52 0.18 0.88 ;
  RECT -0.18 1.22 0.18 1.58 ;
END via8_VX_X3N

VIA via8_VX_X4H DEFAULT
  LAYER M8 ;
  RECT -0.54 -0.58 0.54 0.58 ;
  LAYER TM2 ;
  RECT -0.55 -0.55 0.55 0.55 ;
  LAYER TV2 ;
  RECT -0.53 -0.53 -0.17 -0.17 ;
  RECT -0.53 0.17 -0.17 0.53 ;
  RECT 0.17 -0.53 0.53 -0.17 ;
  RECT 0.17 0.17 0.53 0.53 ;
END via8_VX_X4H

VIA via8_VX_X4E DEFAULT
  LAYER M8 ;
  RECT -0.19 -0.58 0.89 0.58 ;
  LAYER TM2 ;
  RECT -0.2 -0.55 0.9 0.55 ;
  LAYER TV2 ;
  RECT -0.18 -0.53 0.18 -0.17 ;
  RECT -0.18 0.17 0.18 0.53 ;
  RECT 0.52 -0.53 0.88 -0.17 ;
  RECT 0.52 0.17 0.88 0.53 ;
END via8_VX_X4E

VIA via8_VX_X4W DEFAULT
  LAYER M8 ;
  RECT -0.89 -0.58 0.19 0.58 ;
  LAYER TM2 ;
  RECT -0.9 -0.55 0.2 0.55 ;
  LAYER TV2 ;
  RECT -0.88 -0.53 -0.52 -0.17 ;
  RECT -0.88 0.17 -0.52 0.53 ;
  RECT -0.18 -0.53 0.18 -0.17 ;
  RECT -0.18 0.17 0.18 0.53 ;
END via8_VX_X4W

VIA via8_VX_X4S DEFAULT
  LAYER M8 ;
  RECT -0.54 -0.93 0.54 0.23 ;
  LAYER TM2 ;
  RECT -0.55 -0.9 0.55 0.2 ;
  LAYER TV2 ;
  RECT -0.53 -0.88 -0.17 -0.52 ;
  RECT -0.53 -0.18 -0.17 0.18 ;
  RECT 0.17 -0.88 0.53 -0.52 ;
  RECT 0.17 -0.18 0.53 0.18 ;
END via8_VX_X4S

VIA via8_VX_X4N DEFAULT
  LAYER M8 ;
  RECT -0.54 -0.23 0.54 0.93 ;
  LAYER TM2 ;
  RECT -0.55 -0.2 0.55 0.9 ;
  LAYER TV2 ;
  RECT -0.53 -0.18 -0.17 0.18 ;
  RECT -0.53 0.52 -0.17 0.88 ;
  RECT 0.17 -0.18 0.53 0.18 ;
  RECT 0.17 0.52 0.53 0.88 ;
END via8_VX_X4N

VIA via9_RDV_X2H DEFAULT
  LAYER TM2 ;
  RECT -5.5 -2.5 5.5 2.5 ;
  LAYER RDL ;
  RECT -6 -3 6 3 ;
  LAYER RDV ;
  RECT -4.5 -1.5 -1.5 1.5 ;
  RECT 1.5 -1.5 4.5 1.5 ;
END via9_RDV_X2H

VIA via9_RDV_X2E DEFAULT
  LAYER TM2 ;
  RECT -2.5 -2.5 8.5 2.5 ;
  LAYER RDL ;
  RECT -3 -3 9 3 ;
  LAYER RDV ;
  RECT -1.5 -1.5 1.5 1.5 ;
  RECT 4.5 -1.5 7.5 1.5 ;
END via9_RDV_X2E

VIA via9_RDV_X2W DEFAULT
  LAYER TM2 ;
  RECT -8.5 -2.5 2.5 2.5 ;
  LAYER RDL ;
  RECT -9 -3 3 3 ;
  LAYER RDV ;
  RECT -7.5 -1.5 -4.5 1.5 ;
  RECT -1.5 -1.5 1.5 1.5 ;
END via9_RDV_X2W

VIA via9_RDV_X2V DEFAULT
  LAYER TM2 ;
  RECT -2.5 -5.5 2.5 5.5 ;
  LAYER RDL ;
  RECT -3 -6 3 6 ;
  LAYER RDV ;
  RECT -1.5 -4.5 1.5 -1.5 ;
  RECT -1.5 1.5 1.5 4.5 ;
END via9_RDV_X2V

VIA via9_RDV_X2S DEFAULT
  LAYER TM2 ;
  RECT -2.5 -8.5 2.5 2.5 ;
  LAYER RDL ;
  RECT -3 -9 3 3 ;
  LAYER RDV ;
  RECT -1.5 -7.5 1.5 -4.5 ;
  RECT -1.5 -1.5 1.5 1.5 ;
END via9_RDV_X2S

VIA via9_RDV_X2N DEFAULT
  LAYER TM2 ;
  RECT -2.5 -2.5 2.5 8.5 ;
  LAYER RDL ;
  RECT -3 -3 3 9 ;
  LAYER RDV ;
  RECT -1.5 -1.5 1.5 1.5 ;
  RECT -1.5 4.5 1.5 7.5 ;
END via9_RDV_X2N

VIA via9_RDV_X3H DEFAULT
  LAYER TM2 ;
  RECT -8.5 -2.5 8.5 2.5 ;
  LAYER RDL ;
  RECT -9 -3 9 3 ;
  LAYER RDV ;
  RECT -7.5 -1.5 -4.5 1.5 ;
  RECT -1.5 -1.5 1.5 1.5 ;
  RECT 4.5 -1.5 7.5 1.5 ;
END via9_RDV_X3H

VIA via9_RDV_X3E DEFAULT
  LAYER TM2 ;
  RECT -2.5 -2.5 14.5 2.5 ;
  LAYER RDL ;
  RECT -3 -3 15 3 ;
  LAYER RDV ;
  RECT -1.5 -1.5 1.5 1.5 ;
  RECT 4.5 -1.5 7.5 1.5 ;
  RECT 10.5 -1.5 13.5 1.5 ;
END via9_RDV_X3E

VIA via9_RDV_X3W DEFAULT
  LAYER TM2 ;
  RECT -14.5 -2.5 2.5 2.5 ;
  LAYER RDL ;
  RECT -15 -3 3 3 ;
  LAYER RDV ;
  RECT -13.5 -1.5 -10.5 1.5 ;
  RECT -7.5 -1.5 -4.5 1.5 ;
  RECT -1.5 -1.5 1.5 1.5 ;
END via9_RDV_X3W

VIA via9_RDV_X3V DEFAULT
  LAYER TM2 ;
  RECT -2.5 -8.5 2.5 8.5 ;
  LAYER RDL ;
  RECT -3 -9 3 9 ;
  LAYER RDV ;
  RECT -1.5 -7.5 1.5 -4.5 ;
  RECT -1.5 -1.5 1.5 1.5 ;
  RECT -1.5 4.5 1.5 7.5 ;
END via9_RDV_X3V

VIA via9_RDV_X3S DEFAULT
  LAYER TM2 ;
  RECT -2.5 -14.5 2.5 2.5 ;
  LAYER RDL ;
  RECT -3 -15 3 3 ;
  LAYER RDV ;
  RECT -1.5 -13.5 1.5 -10.5 ;
  RECT -1.5 -7.5 1.5 -4.5 ;
  RECT -1.5 -1.5 1.5 1.5 ;
END via9_RDV_X3S

VIA via9_RDV_X3N DEFAULT
  LAYER TM2 ;
  RECT -2.5 -2.5 2.5 14.5 ;
  LAYER RDL ;
  RECT -3 -3 3 15 ;
  LAYER RDV ;
  RECT -1.5 -1.5 1.5 1.5 ;
  RECT -1.5 4.5 1.5 7.5 ;
  RECT -1.5 10.5 1.5 13.5 ;
END via9_RDV_X3N

VIA via9_RDV_X4H DEFAULT
  LAYER TM2 ;
  RECT -5.5 -5.5 5.5 5.5 ;
  LAYER RDL ;
  RECT -6 -6 6 6 ;
  LAYER RDV ;
  RECT -4.5 -4.5 -1.5 -1.5 ;
  RECT -4.5 1.5 -1.5 4.5 ;
  RECT 1.5 -4.5 4.5 -1.5 ;
  RECT 1.5 1.5 4.5 4.5 ;
END via9_RDV_X4H

VIA via9_RDV_X4E DEFAULT
  LAYER TM2 ;
  RECT -2.5 -5.5 8.5 5.5 ;
  LAYER RDL ;
  RECT -3 -6 9 6 ;
  LAYER RDV ;
  RECT -1.5 -4.5 1.5 -1.5 ;
  RECT -1.5 1.5 1.5 4.5 ;
  RECT 4.5 -4.5 7.5 -1.5 ;
  RECT 4.5 1.5 7.5 4.5 ;
END via9_RDV_X4E

VIA via9_RDV_X4W DEFAULT
  LAYER TM2 ;
  RECT -8.5 -5.5 2.5 5.5 ;
  LAYER RDL ;
  RECT -9 -6 3 6 ;
  LAYER RDV ;
  RECT -7.5 -4.5 -4.5 -1.5 ;
  RECT -7.5 1.5 -4.5 4.5 ;
  RECT -1.5 -4.5 1.5 -1.5 ;
  RECT -1.5 1.5 1.5 4.5 ;
END via9_RDV_X4W

VIA via9_RDV_X4S DEFAULT
  LAYER TM2 ;
  RECT -5.5 -8.5 5.5 2.5 ;
  LAYER RDL ;
  RECT -6 -9 6 3 ;
  LAYER RDV ;
  RECT -4.5 -7.5 -1.5 -4.5 ;
  RECT -4.5 -1.5 -1.5 1.5 ;
  RECT 1.5 -7.5 4.5 -4.5 ;
  RECT 1.5 -1.5 4.5 1.5 ;
END via9_RDV_X4S

VIA via9_RDV_X4N DEFAULT
  LAYER TM2 ;
  RECT -5.5 -2.5 5.5 8.5 ;
  LAYER RDL ;
  RECT -6 -3 6 9 ;
  LAYER RDV ;
  RECT -4.5 -1.5 -1.5 1.5 ;
  RECT -4.5 4.5 -1.5 7.5 ;
  RECT 1.5 -1.5 4.5 1.5 ;
  RECT 1.5 4.5 4.5 7.5 ;
END via9_RDV_X4N

VIARULE via1_fat_arr GENERATE
  LAYER M1 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M2 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via1_fat_arr

VIARULE via2_fat_arr GENERATE
  LAYER M2 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M3 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via2_fat_arr

VIARULE via3_fat_arr GENERATE
  LAYER M3 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M4 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via3_fat_arr

VIARULE via4_fat_arr GENERATE
  LAYER M4 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M5 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V4 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via4_fat_arr

VIARULE via5_fat_arr GENERATE
  LAYER M5 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M6 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V5 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via5_fat_arr

VIARULE via6_fat_arr GENERATE
  LAYER M6 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M7 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V6 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via6_fat_arr

VIARULE via7_fat_arr GENERATE
  LAYER M7 ;
  ENCLOSURE 0.03 0.03 ;
  LAYER M8 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER V7 ;
  RECT -0.045 -0.045 0.045 0.045 ;
  SPACING 0.22 BY 0.22 ;
END via7_fat_arr

VIARULE via8_fat_arr GENERATE
  LAYER M8 ;
  ENCLOSURE 0.05 0.05 ;
  LAYER TM2 ;
  ENCLOSURE 0.02 0.02 ;
  LAYER TV2 ;
  RECT -0.18 -0.18 0.18 0.18 ;
  SPACING 0.86 BY 0.86 ;
END via8_fat_arr

END LIBRARY
