* File: rcx_out.net
* Created: Tue Mar 26 09:51:54 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:51:54 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt MAJ3X1  A B C VDD VSS Y
* 
XM11/X1 Y net29 net24 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM8/X1 net24 net13 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM7/X1 Y net14 net23 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM3/X1 net23 net29 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM1/X1 net26 net14 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM2/X1 Y net13 net26 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.8801e-12 PD=2.23088e-05
XM22/X1 Y net14 net25 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.08121e-11 PD=3.35088e-05
XM23/X1 net28 net14 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM24/X1 Y net29 net28 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM0/X1 net25 net13 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM25/X1 Y net13 net27 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM26/X1 net27 net29 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XI3/XM1/X1 net29 C VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9285e-12 PD=1.67888e-05
XI3/XM0/X1 net29 C VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XI2/XM1/X1 net13 A VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9285e-12 PD=1.67888e-05
XI2/XM0/X1 net13 A VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XI0/XM1/X1 net14 B VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=4.9285e-12 PD=1.67888e-05
XI0/XM0/X1 net14 B VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
*
* 
* .include "rcx_out.net.MAJ3X1.pxi"
* BEGIN of "./rcx_out.net.MAJ3X1.pxi"
* File: rcx_out.net.MAJ3X1.pxi
* Created: Tue Mar 26 09:51:54 2019
* 

* END of "./rcx_out.net.MAJ3X1.pxi"
* 
*
.ends
*
*

