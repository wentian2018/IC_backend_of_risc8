* File: rcx_out.net
* Created: Tue Mar 26 09:46:06 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:46:06 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt INVX16  A VDD VSS Y
* 
XM1/X1 Y A VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=8
XM0/X1 Y A VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=8
*
* 
* .include "rcx_out.net.INVX16.pxi"
* BEGIN of "./rcx_out.net.INVX16.pxi"
* File: rcx_out.net.INVX16.pxi
* Created: Tue Mar 26 09:46:06 2019
* 

* END of "./rcx_out.net.INVX16.pxi"
* 
*
.ends
*
*

