* File: rcx_out.net
* Created: Tue Mar 26 09:43:30 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:43:30 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt NOR2X1  A B VDD VSS Y
* 
XM2/X1 Y B net010 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.29593e-11 PD=3.41488e-05
XM1/X1 net010 A VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.29593e-11 PD=3.41488e-05
XM3/X1 Y B VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=5.8465e-12 PD=1.75088e-05
XM0/X1 Y A VSS VSS nch_5_mac_egl4 A=7.4e-07 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=5.276e-13 PS=2.72569e-06
+ AD=5.8465e-12 PD=1.75088e-05
*
* 
* .include "rcx_out.net.NOR2X1.pxi"
* BEGIN of "./rcx_out.net.NOR2X1.pxi"
* File: rcx_out.net.NOR2X1.pxi
* Created: Tue Mar 26 09:43:30 2019
* 

* END of "./rcx_out.net.NOR2X1.pxi"
* 
*
.ends
*
*

