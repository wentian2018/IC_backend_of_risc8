* File: rcx_out.net
* Created: Tue Mar 26 09:51:01 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:51:01 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt OAI21X1  A0 A1 B0 VDD VSS Y
* 
XM11/X1 Y B0 net07 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=7.1147e-12 PD=2.24288e-05
XM0/X1 net07 A1 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=7.0365e-12 PD=2.23888e-05
XM3/X1 net07 A0 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=7.1147e-12 PD=2.24288e-05
XM8/X1 Y B0 VDD VDD pch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=7.1147e-12 PD=2.24288e-05
XM2/X1 net015 A1 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.10805e-11 PD=3.35888e-05
XM1/X1 Y A0 net015 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.12147e-11 PD=3.36288e-05
*
* 
* .include "rcx_out.net.OAI21X1.pxi"
* BEGIN of "./rcx_out.net.OAI21X1.pxi"
* File: rcx_out.net.OAI21X1.pxi
* Created: Tue Mar 26 09:51:01 2019
* 

* END of "./rcx_out.net.OAI21X1.pxi"
* 
*
.ends
*
*

