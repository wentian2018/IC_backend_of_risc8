* File: rcx_out.net
* Created: Tue Mar 26 09:50:07 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* 
* 
* .include "rcx_out.net.pex"
* BEGIN of "./rcx_out.net.pex"
* File: rcx_out.net.pex
* Created: Tue Mar 26 09:50:07 2019
* Program "Calibre xRC"
* Version "v2013.2_35.25"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 

* END of "./rcx_out.net.pex"
* 
.subckt DLYX1  A VDD VSS Y
* 
XM59/X1 net010 net026 net087 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07
+ H=5e-07 NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12
+ PS=5.44569e-06 AD=6.7237e-12 PD=2.22288e-05
XM62/X1 net13 net010 net084 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07
+ H=5e-07 NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12
+ PS=5.44569e-06 AD=6.7237e-12 PD=2.22288e-05
XM60/X1 net087 net026 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM61/X1 net084 net010 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM70/X1 VSS net026 VSS VSS nch_5_mac_egl4 A=3.6e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=3
XM58/X1 net040 A VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM10/X1 net026 A net040 VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=1.49941e-07 HAB=6.59956e-07 AS=1.534e-12 PS=5.44569e-06
+ AD=6.7237e-12 PD=2.22288e-05
XM6/X1 Y net13 VSS VSS nch_5_mac_egl4 A=2.1e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=4
XM72/X1 VSS net13 VSS VSS nch_5_mac_egl4 A=3.6e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=3
XM56/X1 net010 net026 net085 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07
+ H=5e-07 NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12
+ PS=1.08457e-05 AD=1.05437e-11 PD=3.34288e-05
XM39/X1 net085 net026 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM69/X1 VDD net026 VDD VDD pch_5_mac_egl4 A=7.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=3
XM55/X1 net026 A net039 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM19/X1 net039 A VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=1
+ POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM7/X1 Y net13 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07 NF=4
XM71/X1 VDD net13 VDD VDD pch_5_mac_egl4 A=7.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=3
XM48/X1 net083 net010 VDD VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07 H=5e-07
+ NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12 PS=1.08457e-05
+ AD=1.05437e-11 PD=3.34288e-05
XM57/X1 net13 net010 net083 VDD pch_5_mac_egl4 A=4.8e-06 B=7.4e-07 D=1e-07
+ H=5e-07 NF=1 POLYCNN=5e-07 HAT=2.49941e-07 HAB=6.59956e-07 AS=3.532e-12
+ PS=1.08457e-05 AD=1.05437e-11 PD=3.34288e-05
*
* 
* .include "rcx_out.net.DLYX1.pxi"
* BEGIN of "./rcx_out.net.DLYX1.pxi"
* File: rcx_out.net.DLYX1.pxi
* Created: Tue Mar 26 09:50:07 2019
* 

* END of "./rcx_out.net.DLYX1.pxi"
* 
*
.ends
*
*

